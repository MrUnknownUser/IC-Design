// Generator : SpinalHDL v1.12.3    git head : 591e64062329e5e2e2b81f4d52422948053edb97
// Component : AesIterative
// Git hash  : bbee732ce863f54b6bd0cc5b3b23faaf1003bdf0

`timescale 1ns/1ps

module AesIterative (
  input  wire          io_start,
  input  wire          io_decrypt,
  input  wire [127:0]  io_key,
  input  wire [127:0]  io_dataIn,
  output reg  [127:0]  io_dataOut,
  output wire          io_busy,
  output reg           io_done,
  input  wire          clk,
  input  wire          reset
);

  wire       [79:0]   _zz_stateReg_75;
  wire       [39:0]   _zz_stateReg_76;
  wire       [7:0]    _zz_stateReg_77;
  wire       [7:0]    _zz_stateReg_78;
  wire       [7:0]    _zz_stateReg_79;
  wire       [7:0]    _zz_stateReg_80;
  wire       [7:0]    _zz_stateReg_81;
  wire       [7:0]    _zz_stateReg_82;
  wire       [7:0]    _zz_stateReg_83;
  wire       [7:0]    _zz_stateReg_84;
  wire       [7:0]    _zz_stateReg_85;
  wire       [7:0]    _zz_stateReg_86;
  wire       [7:0]    _zz_stateReg_87;
  wire       [7:0]    _zz_stateReg_88;
  wire       [7:0]    _zz_stateReg_89;
  wire       [7:0]    _zz_stateReg_90;
  wire       [7:0]    _zz_stateReg_91;
  reg        [7:0]    _zz__zz_stateReg_4;
  wire       [7:0]    _zz__zz_stateReg_4_1;
  reg        [7:0]    _zz__zz_stateReg_8;
  wire       [7:0]    _zz__zz_stateReg_8_1;
  reg        [7:0]    _zz__zz_stateReg_12;
  wire       [7:0]    _zz__zz_stateReg_12_1;
  reg        [7:0]    _zz__zz_stateReg_16;
  wire       [7:0]    _zz__zz_stateReg_16_1;
  reg        [7:0]    _zz__zz_stateReg_5;
  wire       [7:0]    _zz__zz_stateReg_5_1;
  reg        [7:0]    _zz__zz_stateReg_9;
  wire       [7:0]    _zz__zz_stateReg_9_1;
  reg        [7:0]    _zz__zz_stateReg_13;
  wire       [7:0]    _zz__zz_stateReg_13_1;
  reg        [7:0]    _zz__zz_stateReg_17;
  wire       [7:0]    _zz__zz_stateReg_17_1;
  reg        [7:0]    _zz__zz_stateReg_6;
  wire       [7:0]    _zz__zz_stateReg_6_1;
  reg        [7:0]    _zz__zz_stateReg_10;
  wire       [7:0]    _zz__zz_stateReg_10_1;
  reg        [7:0]    _zz__zz_stateReg_14;
  wire       [7:0]    _zz__zz_stateReg_14_1;
  reg        [7:0]    _zz__zz_stateReg_18;
  wire       [7:0]    _zz__zz_stateReg_18_1;
  reg        [7:0]    _zz__zz_stateReg_7;
  wire       [7:0]    _zz__zz_stateReg_7_1;
  reg        [7:0]    _zz__zz_stateReg_11;
  wire       [7:0]    _zz__zz_stateReg_11_1;
  reg        [7:0]    _zz__zz_stateReg_15;
  wire       [7:0]    _zz__zz_stateReg_15_1;
  reg        [7:0]    _zz__zz_stateReg_19;
  wire       [7:0]    _zz__zz_stateReg_19_1;
  wire       [8:0]    _zz__zz_stateReg_36;
  wire       [8:0]    _zz__zz_stateReg_37;
  wire       [8:0]    _zz__zz_stateReg_38;
  wire       [8:0]    _zz__zz_stateReg_39;
  wire       [8:0]    _zz__zz_stateReg_40;
  wire       [8:0]    _zz__zz_stateReg_41;
  wire       [8:0]    _zz__zz_stateReg_42;
  wire       [8:0]    _zz__zz_stateReg_43;
  wire       [8:0]    _zz__zz_stateReg_44;
  wire       [8:0]    _zz__zz_stateReg_45;
  wire       [8:0]    _zz__zz_stateReg_46;
  wire       [8:0]    _zz__zz_stateReg_47;
  wire       [8:0]    _zz__zz_stateReg_48;
  wire       [8:0]    _zz__zz_stateReg_49;
  wire       [8:0]    _zz__zz_stateReg_50;
  wire       [8:0]    _zz__zz_stateReg_51;
  wire       [8:0]    _zz__zz_stateReg_52;
  wire       [8:0]    _zz__zz_stateReg_53;
  wire       [8:0]    _zz__zz_stateReg_54;
  wire       [8:0]    _zz__zz_stateReg_55;
  wire       [8:0]    _zz__zz_stateReg_56;
  wire       [8:0]    _zz__zz_stateReg_57;
  wire       [8:0]    _zz__zz_stateReg_58;
  wire       [8:0]    _zz__zz_stateReg_59;
  wire       [8:0]    _zz__zz_stateReg_60;
  wire       [8:0]    _zz__zz_stateReg_61;
  wire       [8:0]    _zz__zz_stateReg_62;
  wire       [8:0]    _zz__zz_stateReg_63;
  wire       [8:0]    _zz__zz_stateReg_64;
  wire       [8:0]    _zz__zz_stateReg_65;
  wire       [8:0]    _zz__zz_stateReg_66;
  wire       [8:0]    _zz__zz_stateReg_67;
  wire       [39:0]   _zz__zz_stateReg_68;
  wire       [7:0]    _zz__zz_stateReg_68_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_3;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2_4;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_5;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2_6;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_7;
  wire       [55:0]   _zz__zz_stateReg_69;
  wire       [7:0]    _zz__zz_stateReg_69_1;
  wire       [7:0]    _zz__zz_stateReg_69_2;
  reg        [7:0]    _zz__zz_stateReg_71;
  wire       [7:0]    _zz__zz_stateReg_71_1;
  reg        [7:0]    _zz__zz_stateReg_71_2;
  wire       [7:0]    _zz__zz_stateReg_71_3;
  reg        [7:0]    _zz__zz_stateReg_71_4;
  wire       [7:0]    _zz__zz_stateReg_71_5;
  reg        [7:0]    _zz__zz_stateReg_71_6;
  wire       [7:0]    _zz__zz_stateReg_71_7;
  reg        [7:0]    _zz__zz_stateReg_71_8;
  wire       [55:0]   _zz_stateReg_92;
  wire       [7:0]    _zz_stateReg_93;
  wire       [7:0]    _zz_stateReg_94;
  reg        [7:0]    _zz_invSub_0;
  reg        [7:0]    _zz_invSub_1;
  reg        [7:0]    _zz_invSub_2;
  reg        [7:0]    _zz_invSub_3;
  reg        [7:0]    _zz_invSub_4;
  reg        [7:0]    _zz_invSub_5;
  reg        [7:0]    _zz_invSub_6;
  reg        [7:0]    _zz_invSub_7;
  reg        [7:0]    _zz_invSub_8;
  reg        [7:0]    _zz_invSub_9;
  reg        [7:0]    _zz_invSub_10;
  reg        [7:0]    _zz_invSub_11;
  reg        [7:0]    _zz_invSub_12;
  reg        [7:0]    _zz_invSub_13;
  reg        [7:0]    _zz_invSub_14;
  reg        [7:0]    _zz_invSub_15;
  reg        [7:0]    _zz__zz_roundKeyReg_0_5;
  wire       [7:0]    _zz__zz_roundKeyReg_0_5_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0_5_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_5_3;
  reg        [7:0]    _zz__zz_roundKeyReg_0_5_4;
  wire       [7:0]    _zz__zz_roundKeyReg_0_5_5;
  reg        [7:0]    _zz__zz_roundKeyReg_0_5_6;
  wire       [7:0]    _zz__zz_roundKeyReg_0_5_7;
  wire       [87:0]   _zz__zz_invMixed_0;
  wire       [47:0]   _zz__zz_invMixed_0_1;
  wire       [7:0]    _zz__zz_invMixed_0_2;
  wire       [7:0]    _zz__zz_invMixed_0_3;
  wire       [7:0]    _zz__zz_invMixed_0_4;
  wire       [7:0]    _zz__zz_invMixed_0_5;
  wire       [87:0]   _zz__zz_invMixed_0_6;
  wire       [47:0]   _zz__zz_invMixed_0_7;
  wire       [7:0]    _zz__zz_invMixed_0_8;
  wire       [7:0]    _zz__zz_invMixed_0_9;
  wire       [7:0]    _zz__zz_invMixed_0_10;
  wire       [7:0]    _zz__zz_invMixed_0_11;
  wire       [7:0]    _zz__zz_invMixed_0_12;
  wire       [7:0]    _zz__zz_invMixed_0_13;
  wire       [7:0]    _zz__zz_invMixed_0_14;
  wire       [8:0]    _zz__zz_invMixed_0_5_1;
  wire       [8:0]    _zz__zz_invMixed_0_7_1;
  wire       [8:0]    _zz__zz_invMixed_0_9_1;
  wire       [8:0]    _zz__zz_invMixed_0_10_1;
  wire       [8:0]    _zz__zz_invMixed_0_12_1;
  wire       [8:0]    _zz__zz_invMixed_0_13_1;
  wire       [8:0]    _zz__zz_invMixed_0_14_1;
  wire       [8:0]    _zz__zz_invMixed_0_16;
  wire       [8:0]    _zz__zz_invMixed_0_18;
  wire       [8:0]    _zz__zz_invMixed_0_19;
  wire       [8:0]    _zz__zz_invMixed_0_20;
  wire       [8:0]    _zz__zz_invMixed_0_22;
  wire       [8:0]    _zz__zz_invMixed_0_24;
  wire       [8:0]    _zz__zz_invMixed_0_25;
  wire       [8:0]    _zz__zz_invMixed_0_27;
  wire       [8:0]    _zz__zz_invMixed_0_28;
  wire       [8:0]    _zz__zz_invMixed_0_30;
  wire       [8:0]    _zz__zz_invMixed_0_32;
  wire       [8:0]    _zz__zz_invMixed_1;
  wire       [8:0]    _zz__zz_invMixed_1_2;
  wire       [8:0]    _zz__zz_invMixed_1_4;
  wire       [8:0]    _zz__zz_invMixed_1_5;
  wire       [8:0]    _zz__zz_invMixed_1_7;
  wire       [8:0]    _zz__zz_invMixed_1_9;
  wire       [8:0]    _zz__zz_invMixed_1_10;
  wire       [8:0]    _zz__zz_invMixed_1_12;
  wire       [8:0]    _zz__zz_invMixed_1_13;
  wire       [8:0]    _zz__zz_invMixed_1_14;
  wire       [8:0]    _zz__zz_invMixed_1_16;
  wire       [8:0]    _zz__zz_invMixed_1_18;
  wire       [8:0]    _zz__zz_invMixed_1_19;
  wire       [8:0]    _zz__zz_invMixed_1_20;
  wire       [8:0]    _zz__zz_invMixed_1_22;
  wire       [8:0]    _zz__zz_invMixed_1_24;
  wire       [8:0]    _zz__zz_invMixed_1_25;
  wire       [8:0]    _zz__zz_invMixed_1_27;
  wire       [8:0]    _zz__zz_invMixed_2;
  wire       [8:0]    _zz__zz_invMixed_2_2;
  wire       [8:0]    _zz__zz_invMixed_2_4;
  wire       [8:0]    _zz__zz_invMixed_2_5;
  wire       [8:0]    _zz__zz_invMixed_2_7;
  wire       [8:0]    _zz__zz_invMixed_2_8;
  wire       [8:0]    _zz__zz_invMixed_2_10;
  wire       [8:0]    _zz__zz_invMixed_2_12;
  wire       [8:0]    _zz__zz_invMixed_2_13;
  wire       [8:0]    _zz__zz_invMixed_2_15;
  wire       [8:0]    _zz__zz_invMixed_2_17;
  wire       [8:0]    _zz__zz_invMixed_2_18;
  wire       [8:0]    _zz__zz_invMixed_2_20;
  wire       [8:0]    _zz__zz_invMixed_2_21;
  wire       [8:0]    _zz__zz_invMixed_2_22;
  wire       [8:0]    _zz__zz_invMixed_2_24;
  wire       [8:0]    _zz__zz_invMixed_2_26;
  wire       [8:0]    _zz__zz_invMixed_2_27;
  wire       [8:0]    _zz__zz_invMixed_3;
  wire       [8:0]    _zz__zz_invMixed_3_2;
  wire       [8:0]    _zz__zz_invMixed_3_4;
  wire       [8:0]    _zz__zz_invMixed_3_5;
  wire       [8:0]    _zz__zz_invMixed_3_6;
  wire       [8:0]    _zz__zz_invMixed_3_8;
  wire       [8:0]    _zz__zz_invMixed_3_10;
  wire       [8:0]    _zz__zz_invMixed_3_11;
  wire       [8:0]    _zz__zz_invMixed_3_13;
  wire       [8:0]    _zz__zz_invMixed_3_14;
  wire       [8:0]    _zz__zz_invMixed_3_16;
  wire       [8:0]    _zz__zz_invMixed_3_18;
  wire       [8:0]    _zz__zz_invMixed_3_19;
  wire       [8:0]    _zz__zz_invMixed_3_21;
  wire       [8:0]    _zz__zz_invMixed_3_23;
  wire       [8:0]    _zz__zz_invMixed_3_24;
  wire       [8:0]    _zz__zz_invMixed_3_26;
  wire       [8:0]    _zz__zz_invMixed_3_27;
  wire       [7:0]    _zz_invMixed_0_33;
  wire       [7:0]    _zz_invMixed_0_34;
  wire                _zz_invMixed_0_35;
  wire       [7:0]    _zz_invMixed_0_36;
  wire       [7:0]    _zz_invMixed_0_37;
  wire       [7:0]    _zz_invMixed_0_38;
  wire                _zz_invMixed_0_39;
  wire       [7:0]    _zz_invMixed_0_40;
  wire                _zz_invMixed_0_41;
  wire       [7:0]    _zz_invMixed_0_42;
  wire                _zz_invMixed_1_28;
  wire       [7:0]    _zz_invMixed_1_29;
  wire       [7:0]    _zz_invMixed_1_30;
  wire       [7:0]    _zz_invMixed_1_31;
  wire                _zz_invMixed_1_32;
  wire       [7:0]    _zz_invMixed_1_33;
  wire                _zz_invMixed_1_34;
  wire       [7:0]    _zz_invMixed_1_35;
  wire                _zz_invMixed_1_36;
  wire       [7:0]    _zz_invMixed_1_37;
  wire       [7:0]    _zz_invMixed_1_38;
  wire       [7:0]    _zz_invMixed_1_39;
  wire       [7:0]    _zz_invMixed_2_28;
  wire       [7:0]    _zz_invMixed_2_29;
  wire                _zz_invMixed_2_30;
  wire       [7:0]    _zz_invMixed_2_31;
  wire                _zz_invMixed_2_32;
  wire       [7:0]    _zz_invMixed_2_33;
  wire                _zz_invMixed_2_34;
  wire       [7:0]    _zz_invMixed_2_35;
  wire       [7:0]    _zz_invMixed_2_36;
  wire       [7:0]    _zz_invMixed_2_37;
  wire       [7:0]    _zz_invMixed_2_38;
  wire       [7:0]    _zz_invMixed_3_28;
  wire       [7:0]    _zz_invMixed_3_29;
  wire       [7:0]    _zz_invMixed_3_30;
  wire       [7:0]    _zz_invMixed_3_31;
  wire       [7:0]    _zz_invMixed_3_32;
  wire       [7:0]    _zz_invMixed_3_33;
  wire       [7:0]    _zz_invMixed_3_34;
  wire       [8:0]    _zz__zz_invMixed_4_4;
  wire       [8:0]    _zz__zz_invMixed_4_6;
  wire       [8:0]    _zz__zz_invMixed_4_8;
  wire       [8:0]    _zz__zz_invMixed_4_9;
  wire       [8:0]    _zz__zz_invMixed_4_11;
  wire       [8:0]    _zz__zz_invMixed_4_12;
  wire       [8:0]    _zz__zz_invMixed_4_13;
  wire       [8:0]    _zz__zz_invMixed_4_15;
  wire       [8:0]    _zz__zz_invMixed_4_17;
  wire       [8:0]    _zz__zz_invMixed_4_18;
  wire       [8:0]    _zz__zz_invMixed_4_19;
  wire       [8:0]    _zz__zz_invMixed_4_21;
  wire       [8:0]    _zz__zz_invMixed_4_23;
  wire       [8:0]    _zz__zz_invMixed_4_24;
  wire       [8:0]    _zz__zz_invMixed_4_26;
  wire       [8:0]    _zz__zz_invMixed_4_27;
  wire       [8:0]    _zz__zz_invMixed_4_29;
  wire       [8:0]    _zz__zz_invMixed_4_31;
  wire       [8:0]    _zz__zz_invMixed_5;
  wire       [8:0]    _zz__zz_invMixed_5_2;
  wire       [8:0]    _zz__zz_invMixed_5_4;
  wire       [8:0]    _zz__zz_invMixed_5_5;
  wire       [8:0]    _zz__zz_invMixed_5_7;
  wire       [8:0]    _zz__zz_invMixed_5_9;
  wire       [8:0]    _zz__zz_invMixed_5_10;
  wire       [8:0]    _zz__zz_invMixed_5_12;
  wire       [8:0]    _zz__zz_invMixed_5_13;
  wire       [8:0]    _zz__zz_invMixed_5_14;
  wire       [8:0]    _zz__zz_invMixed_5_16;
  wire       [8:0]    _zz__zz_invMixed_5_18;
  wire       [8:0]    _zz__zz_invMixed_5_19;
  wire       [8:0]    _zz__zz_invMixed_5_20;
  wire       [8:0]    _zz__zz_invMixed_5_22;
  wire       [8:0]    _zz__zz_invMixed_5_24;
  wire       [8:0]    _zz__zz_invMixed_5_25;
  wire       [8:0]    _zz__zz_invMixed_5_27;
  wire       [8:0]    _zz__zz_invMixed_6;
  wire       [8:0]    _zz__zz_invMixed_6_2;
  wire       [8:0]    _zz__zz_invMixed_6_4;
  wire       [8:0]    _zz__zz_invMixed_6_5;
  wire       [8:0]    _zz__zz_invMixed_6_7;
  wire       [8:0]    _zz__zz_invMixed_6_8;
  wire       [8:0]    _zz__zz_invMixed_6_10;
  wire       [8:0]    _zz__zz_invMixed_6_12;
  wire       [8:0]    _zz__zz_invMixed_6_13;
  wire       [8:0]    _zz__zz_invMixed_6_15;
  wire       [8:0]    _zz__zz_invMixed_6_17;
  wire       [8:0]    _zz__zz_invMixed_6_18;
  wire       [8:0]    _zz__zz_invMixed_6_20;
  wire       [8:0]    _zz__zz_invMixed_6_21;
  wire       [8:0]    _zz__zz_invMixed_6_22;
  wire       [8:0]    _zz__zz_invMixed_6_24;
  wire       [8:0]    _zz__zz_invMixed_6_26;
  wire       [8:0]    _zz__zz_invMixed_6_27;
  wire       [8:0]    _zz__zz_invMixed_7;
  wire       [8:0]    _zz__zz_invMixed_7_2;
  wire       [8:0]    _zz__zz_invMixed_7_4;
  wire       [8:0]    _zz__zz_invMixed_7_5;
  wire       [8:0]    _zz__zz_invMixed_7_6;
  wire       [8:0]    _zz__zz_invMixed_7_8;
  wire       [8:0]    _zz__zz_invMixed_7_10;
  wire       [8:0]    _zz__zz_invMixed_7_11;
  wire       [8:0]    _zz__zz_invMixed_7_13;
  wire       [8:0]    _zz__zz_invMixed_7_14;
  wire       [8:0]    _zz__zz_invMixed_7_16;
  wire       [8:0]    _zz__zz_invMixed_7_18;
  wire       [8:0]    _zz__zz_invMixed_7_19;
  wire       [8:0]    _zz__zz_invMixed_7_21;
  wire       [8:0]    _zz__zz_invMixed_7_23;
  wire       [8:0]    _zz__zz_invMixed_7_24;
  wire       [8:0]    _zz__zz_invMixed_7_26;
  wire       [8:0]    _zz__zz_invMixed_7_27;
  wire       [7:0]    _zz_invMixed_4_32;
  wire       [7:0]    _zz_invMixed_4_33;
  wire                _zz_invMixed_4_34;
  wire       [7:0]    _zz_invMixed_4_35;
  wire       [7:0]    _zz_invMixed_4_36;
  wire       [7:0]    _zz_invMixed_4_37;
  wire                _zz_invMixed_4_38;
  wire       [7:0]    _zz_invMixed_4_39;
  wire                _zz_invMixed_4_40;
  wire       [7:0]    _zz_invMixed_4_41;
  wire                _zz_invMixed_5_28;
  wire       [7:0]    _zz_invMixed_5_29;
  wire       [7:0]    _zz_invMixed_5_30;
  wire       [7:0]    _zz_invMixed_5_31;
  wire                _zz_invMixed_5_32;
  wire       [7:0]    _zz_invMixed_5_33;
  wire                _zz_invMixed_5_34;
  wire       [7:0]    _zz_invMixed_5_35;
  wire                _zz_invMixed_5_36;
  wire       [7:0]    _zz_invMixed_5_37;
  wire       [7:0]    _zz_invMixed_5_38;
  wire       [7:0]    _zz_invMixed_5_39;
  wire       [7:0]    _zz_invMixed_6_28;
  wire       [7:0]    _zz_invMixed_6_29;
  wire                _zz_invMixed_6_30;
  wire       [7:0]    _zz_invMixed_6_31;
  wire                _zz_invMixed_6_32;
  wire       [7:0]    _zz_invMixed_6_33;
  wire                _zz_invMixed_6_34;
  wire       [7:0]    _zz_invMixed_6_35;
  wire       [7:0]    _zz_invMixed_6_36;
  wire       [7:0]    _zz_invMixed_6_37;
  wire       [7:0]    _zz_invMixed_6_38;
  wire       [7:0]    _zz_invMixed_7_28;
  wire       [7:0]    _zz_invMixed_7_29;
  wire       [7:0]    _zz_invMixed_7_30;
  wire       [7:0]    _zz_invMixed_7_31;
  wire       [7:0]    _zz_invMixed_7_32;
  wire       [7:0]    _zz_invMixed_7_33;
  wire       [7:0]    _zz_invMixed_7_34;
  wire       [8:0]    _zz__zz_invMixed_8_4;
  wire       [8:0]    _zz__zz_invMixed_8_6;
  wire       [8:0]    _zz__zz_invMixed_8_8;
  wire       [8:0]    _zz__zz_invMixed_8_9;
  wire       [8:0]    _zz__zz_invMixed_8_11;
  wire       [8:0]    _zz__zz_invMixed_8_12;
  wire       [8:0]    _zz__zz_invMixed_8_13;
  wire       [8:0]    _zz__zz_invMixed_8_15;
  wire       [8:0]    _zz__zz_invMixed_8_17;
  wire       [8:0]    _zz__zz_invMixed_8_18;
  wire       [8:0]    _zz__zz_invMixed_8_19;
  wire       [8:0]    _zz__zz_invMixed_8_21;
  wire       [8:0]    _zz__zz_invMixed_8_23;
  wire       [8:0]    _zz__zz_invMixed_8_24;
  wire       [8:0]    _zz__zz_invMixed_8_26;
  wire       [8:0]    _zz__zz_invMixed_8_27;
  wire       [8:0]    _zz__zz_invMixed_8_29;
  wire       [8:0]    _zz__zz_invMixed_8_31;
  wire       [8:0]    _zz__zz_invMixed_9;
  wire       [8:0]    _zz__zz_invMixed_9_2;
  wire       [8:0]    _zz__zz_invMixed_9_4;
  wire       [8:0]    _zz__zz_invMixed_9_5;
  wire       [8:0]    _zz__zz_invMixed_9_7;
  wire       [8:0]    _zz__zz_invMixed_9_9;
  wire       [8:0]    _zz__zz_invMixed_9_10;
  wire       [8:0]    _zz__zz_invMixed_9_12;
  wire       [8:0]    _zz__zz_invMixed_9_13;
  wire       [8:0]    _zz__zz_invMixed_9_14;
  wire       [8:0]    _zz__zz_invMixed_9_16;
  wire       [8:0]    _zz__zz_invMixed_9_18;
  wire       [8:0]    _zz__zz_invMixed_9_19;
  wire       [8:0]    _zz__zz_invMixed_9_20;
  wire       [8:0]    _zz__zz_invMixed_9_22;
  wire       [8:0]    _zz__zz_invMixed_9_24;
  wire       [8:0]    _zz__zz_invMixed_9_25;
  wire       [8:0]    _zz__zz_invMixed_9_27;
  wire       [8:0]    _zz__zz_invMixed_10;
  wire       [8:0]    _zz__zz_invMixed_10_2;
  wire       [8:0]    _zz__zz_invMixed_10_4;
  wire       [8:0]    _zz__zz_invMixed_10_5;
  wire       [8:0]    _zz__zz_invMixed_10_7;
  wire       [8:0]    _zz__zz_invMixed_10_8;
  wire       [8:0]    _zz__zz_invMixed_10_10;
  wire       [8:0]    _zz__zz_invMixed_10_12;
  wire       [8:0]    _zz__zz_invMixed_10_13;
  wire       [8:0]    _zz__zz_invMixed_10_15;
  wire       [8:0]    _zz__zz_invMixed_10_17;
  wire       [8:0]    _zz__zz_invMixed_10_18;
  wire       [8:0]    _zz__zz_invMixed_10_20;
  wire       [8:0]    _zz__zz_invMixed_10_21;
  wire       [8:0]    _zz__zz_invMixed_10_22;
  wire       [8:0]    _zz__zz_invMixed_10_24;
  wire       [8:0]    _zz__zz_invMixed_10_26;
  wire       [8:0]    _zz__zz_invMixed_10_27;
  wire       [8:0]    _zz__zz_invMixed_11;
  wire       [8:0]    _zz__zz_invMixed_11_2;
  wire       [8:0]    _zz__zz_invMixed_11_4;
  wire       [8:0]    _zz__zz_invMixed_11_5;
  wire       [8:0]    _zz__zz_invMixed_11_6;
  wire       [8:0]    _zz__zz_invMixed_11_8;
  wire       [8:0]    _zz__zz_invMixed_11_10;
  wire       [8:0]    _zz__zz_invMixed_11_11;
  wire       [8:0]    _zz__zz_invMixed_11_13;
  wire       [8:0]    _zz__zz_invMixed_11_14;
  wire       [8:0]    _zz__zz_invMixed_11_16;
  wire       [8:0]    _zz__zz_invMixed_11_18;
  wire       [8:0]    _zz__zz_invMixed_11_19;
  wire       [8:0]    _zz__zz_invMixed_11_21;
  wire       [8:0]    _zz__zz_invMixed_11_23;
  wire       [8:0]    _zz__zz_invMixed_11_24;
  wire       [8:0]    _zz__zz_invMixed_11_26;
  wire       [8:0]    _zz__zz_invMixed_11_27;
  wire       [7:0]    _zz_invMixed_8_32;
  wire       [7:0]    _zz_invMixed_8_33;
  wire                _zz_invMixed_8_34;
  wire       [7:0]    _zz_invMixed_8_35;
  wire       [7:0]    _zz_invMixed_8_36;
  wire       [7:0]    _zz_invMixed_8_37;
  wire                _zz_invMixed_8_38;
  wire       [7:0]    _zz_invMixed_8_39;
  wire                _zz_invMixed_8_40;
  wire       [7:0]    _zz_invMixed_8_41;
  wire                _zz_invMixed_9_28;
  wire       [7:0]    _zz_invMixed_9_29;
  wire       [7:0]    _zz_invMixed_9_30;
  wire       [7:0]    _zz_invMixed_9_31;
  wire                _zz_invMixed_9_32;
  wire       [7:0]    _zz_invMixed_9_33;
  wire                _zz_invMixed_9_34;
  wire       [7:0]    _zz_invMixed_9_35;
  wire                _zz_invMixed_9_36;
  wire       [7:0]    _zz_invMixed_9_37;
  wire       [7:0]    _zz_invMixed_9_38;
  wire       [7:0]    _zz_invMixed_9_39;
  wire       [7:0]    _zz_invMixed_10_28;
  wire       [7:0]    _zz_invMixed_10_29;
  wire                _zz_invMixed_10_30;
  wire       [7:0]    _zz_invMixed_10_31;
  wire                _zz_invMixed_10_32;
  wire       [7:0]    _zz_invMixed_10_33;
  wire                _zz_invMixed_10_34;
  wire       [7:0]    _zz_invMixed_10_35;
  wire       [7:0]    _zz_invMixed_10_36;
  wire       [7:0]    _zz_invMixed_10_37;
  wire       [7:0]    _zz_invMixed_10_38;
  wire       [7:0]    _zz_invMixed_11_28;
  wire       [7:0]    _zz_invMixed_11_29;
  wire       [7:0]    _zz_invMixed_11_30;
  wire       [7:0]    _zz_invMixed_11_31;
  wire       [7:0]    _zz_invMixed_11_32;
  wire       [7:0]    _zz_invMixed_11_33;
  wire       [7:0]    _zz_invMixed_11_34;
  wire       [8:0]    _zz__zz_invMixed_12_4;
  wire       [8:0]    _zz__zz_invMixed_12_6;
  wire       [8:0]    _zz__zz_invMixed_12_8;
  wire       [8:0]    _zz__zz_invMixed_12_9;
  wire       [8:0]    _zz__zz_invMixed_12_11;
  wire       [8:0]    _zz__zz_invMixed_12_12;
  wire       [8:0]    _zz__zz_invMixed_12_13;
  wire       [8:0]    _zz__zz_invMixed_12_15;
  wire       [8:0]    _zz__zz_invMixed_12_17;
  wire       [8:0]    _zz__zz_invMixed_12_18;
  wire       [8:0]    _zz__zz_invMixed_12_19;
  wire       [8:0]    _zz__zz_invMixed_12_21;
  wire       [8:0]    _zz__zz_invMixed_12_23;
  wire       [8:0]    _zz__zz_invMixed_12_24;
  wire       [8:0]    _zz__zz_invMixed_12_26;
  wire       [8:0]    _zz__zz_invMixed_12_27;
  wire       [8:0]    _zz__zz_invMixed_12_29;
  wire       [8:0]    _zz__zz_invMixed_12_31;
  wire       [8:0]    _zz__zz_invMixed_13;
  wire       [8:0]    _zz__zz_invMixed_13_2;
  wire       [8:0]    _zz__zz_invMixed_13_4;
  wire       [8:0]    _zz__zz_invMixed_13_5;
  wire       [8:0]    _zz__zz_invMixed_13_7;
  wire       [8:0]    _zz__zz_invMixed_13_9;
  wire       [8:0]    _zz__zz_invMixed_13_10;
  wire       [8:0]    _zz__zz_invMixed_13_12;
  wire       [8:0]    _zz__zz_invMixed_13_13;
  wire       [8:0]    _zz__zz_invMixed_13_14;
  wire       [8:0]    _zz__zz_invMixed_13_16;
  wire       [8:0]    _zz__zz_invMixed_13_18;
  wire       [8:0]    _zz__zz_invMixed_13_19;
  wire       [8:0]    _zz__zz_invMixed_13_20;
  wire       [8:0]    _zz__zz_invMixed_13_22;
  wire       [8:0]    _zz__zz_invMixed_13_24;
  wire       [8:0]    _zz__zz_invMixed_13_25;
  wire       [8:0]    _zz__zz_invMixed_13_27;
  wire       [8:0]    _zz__zz_invMixed_14;
  wire       [8:0]    _zz__zz_invMixed_14_2;
  wire       [8:0]    _zz__zz_invMixed_14_4;
  wire       [8:0]    _zz__zz_invMixed_14_5;
  wire       [8:0]    _zz__zz_invMixed_14_7;
  wire       [8:0]    _zz__zz_invMixed_14_8;
  wire       [8:0]    _zz__zz_invMixed_14_10;
  wire       [8:0]    _zz__zz_invMixed_14_12;
  wire       [8:0]    _zz__zz_invMixed_14_13;
  wire       [8:0]    _zz__zz_invMixed_14_15;
  wire       [8:0]    _zz__zz_invMixed_14_17;
  wire       [8:0]    _zz__zz_invMixed_14_18;
  wire       [8:0]    _zz__zz_invMixed_14_20;
  wire       [8:0]    _zz__zz_invMixed_14_21;
  wire       [8:0]    _zz__zz_invMixed_14_22;
  wire       [8:0]    _zz__zz_invMixed_14_24;
  wire       [8:0]    _zz__zz_invMixed_14_26;
  wire       [8:0]    _zz__zz_invMixed_14_27;
  wire       [8:0]    _zz__zz_invMixed_15;
  wire       [8:0]    _zz__zz_invMixed_15_2;
  wire       [8:0]    _zz__zz_invMixed_15_4;
  wire       [8:0]    _zz__zz_invMixed_15_5;
  wire       [8:0]    _zz__zz_invMixed_15_6;
  wire       [8:0]    _zz__zz_invMixed_15_8;
  wire       [8:0]    _zz__zz_invMixed_15_10;
  wire       [8:0]    _zz__zz_invMixed_15_11;
  wire       [8:0]    _zz__zz_invMixed_15_13;
  wire       [8:0]    _zz__zz_invMixed_15_14;
  wire       [8:0]    _zz__zz_invMixed_15_16;
  wire       [8:0]    _zz__zz_invMixed_15_18;
  wire       [8:0]    _zz__zz_invMixed_15_19;
  wire       [8:0]    _zz__zz_invMixed_15_21;
  wire       [8:0]    _zz__zz_invMixed_15_23;
  wire       [8:0]    _zz__zz_invMixed_15_24;
  wire       [8:0]    _zz__zz_invMixed_15_26;
  wire       [8:0]    _zz__zz_invMixed_15_27;
  wire       [7:0]    _zz_invMixed_12_32;
  wire       [7:0]    _zz_invMixed_12_33;
  wire                _zz_invMixed_12_34;
  wire       [7:0]    _zz_invMixed_12_35;
  wire       [7:0]    _zz_invMixed_12_36;
  wire       [7:0]    _zz_invMixed_12_37;
  wire                _zz_invMixed_12_38;
  wire       [7:0]    _zz_invMixed_12_39;
  wire                _zz_invMixed_12_40;
  wire       [7:0]    _zz_invMixed_12_41;
  wire                _zz_invMixed_13_28;
  wire       [7:0]    _zz_invMixed_13_29;
  wire       [7:0]    _zz_invMixed_13_30;
  wire       [7:0]    _zz_invMixed_13_31;
  wire                _zz_invMixed_13_32;
  wire       [7:0]    _zz_invMixed_13_33;
  wire                _zz_invMixed_13_34;
  wire       [7:0]    _zz_invMixed_13_35;
  wire                _zz_invMixed_13_36;
  wire       [7:0]    _zz_invMixed_13_37;
  wire       [7:0]    _zz_invMixed_13_38;
  wire       [7:0]    _zz_invMixed_13_39;
  wire       [7:0]    _zz_invMixed_14_28;
  wire       [7:0]    _zz_invMixed_14_29;
  wire                _zz_invMixed_14_30;
  wire       [7:0]    _zz_invMixed_14_31;
  wire                _zz_invMixed_14_32;
  wire       [7:0]    _zz_invMixed_14_33;
  wire                _zz_invMixed_14_34;
  wire       [7:0]    _zz_invMixed_14_35;
  wire       [7:0]    _zz_invMixed_14_36;
  wire       [7:0]    _zz_invMixed_14_37;
  wire       [7:0]    _zz_invMixed_14_38;
  wire       [7:0]    _zz_invMixed_15_28;
  wire       [7:0]    _zz_invMixed_15_29;
  wire       [7:0]    _zz_invMixed_15_30;
  wire       [7:0]    _zz_invMixed_15_31;
  wire       [7:0]    _zz_invMixed_15_32;
  wire       [7:0]    _zz_invMixed_15_33;
  wire       [7:0]    _zz_invMixed_15_34;
  wire       [39:0]   _zz_stateReg_95;
  wire       [7:0]    _zz_stateReg_96;
  wire       [7:0]    sboxRom_0;
  wire       [7:0]    sboxRom_1;
  wire       [7:0]    sboxRom_2;
  wire       [7:0]    sboxRom_3;
  wire       [7:0]    sboxRom_4;
  wire       [7:0]    sboxRom_5;
  wire       [7:0]    sboxRom_6;
  wire       [7:0]    sboxRom_7;
  wire       [7:0]    sboxRom_8;
  wire       [7:0]    sboxRom_9;
  wire       [7:0]    sboxRom_10;
  wire       [7:0]    sboxRom_11;
  wire       [7:0]    sboxRom_12;
  wire       [7:0]    sboxRom_13;
  wire       [7:0]    sboxRom_14;
  wire       [7:0]    sboxRom_15;
  wire       [7:0]    sboxRom_16;
  wire       [7:0]    sboxRom_17;
  wire       [7:0]    sboxRom_18;
  wire       [7:0]    sboxRom_19;
  wire       [7:0]    sboxRom_20;
  wire       [7:0]    sboxRom_21;
  wire       [7:0]    sboxRom_22;
  wire       [7:0]    sboxRom_23;
  wire       [7:0]    sboxRom_24;
  wire       [7:0]    sboxRom_25;
  wire       [7:0]    sboxRom_26;
  wire       [7:0]    sboxRom_27;
  wire       [7:0]    sboxRom_28;
  wire       [7:0]    sboxRom_29;
  wire       [7:0]    sboxRom_30;
  wire       [7:0]    sboxRom_31;
  wire       [7:0]    sboxRom_32;
  wire       [7:0]    sboxRom_33;
  wire       [7:0]    sboxRom_34;
  wire       [7:0]    sboxRom_35;
  wire       [7:0]    sboxRom_36;
  wire       [7:0]    sboxRom_37;
  wire       [7:0]    sboxRom_38;
  wire       [7:0]    sboxRom_39;
  wire       [7:0]    sboxRom_40;
  wire       [7:0]    sboxRom_41;
  wire       [7:0]    sboxRom_42;
  wire       [7:0]    sboxRom_43;
  wire       [7:0]    sboxRom_44;
  wire       [7:0]    sboxRom_45;
  wire       [7:0]    sboxRom_46;
  wire       [7:0]    sboxRom_47;
  wire       [7:0]    sboxRom_48;
  wire       [7:0]    sboxRom_49;
  wire       [7:0]    sboxRom_50;
  wire       [7:0]    sboxRom_51;
  wire       [7:0]    sboxRom_52;
  wire       [7:0]    sboxRom_53;
  wire       [7:0]    sboxRom_54;
  wire       [7:0]    sboxRom_55;
  wire       [7:0]    sboxRom_56;
  wire       [7:0]    sboxRom_57;
  wire       [7:0]    sboxRom_58;
  wire       [7:0]    sboxRom_59;
  wire       [7:0]    sboxRom_60;
  wire       [7:0]    sboxRom_61;
  wire       [7:0]    sboxRom_62;
  wire       [7:0]    sboxRom_63;
  wire       [7:0]    sboxRom_64;
  wire       [7:0]    sboxRom_65;
  wire       [7:0]    sboxRom_66;
  wire       [7:0]    sboxRom_67;
  wire       [7:0]    sboxRom_68;
  wire       [7:0]    sboxRom_69;
  wire       [7:0]    sboxRom_70;
  wire       [7:0]    sboxRom_71;
  wire       [7:0]    sboxRom_72;
  wire       [7:0]    sboxRom_73;
  wire       [7:0]    sboxRom_74;
  wire       [7:0]    sboxRom_75;
  wire       [7:0]    sboxRom_76;
  wire       [7:0]    sboxRom_77;
  wire       [7:0]    sboxRom_78;
  wire       [7:0]    sboxRom_79;
  wire       [7:0]    sboxRom_80;
  wire       [7:0]    sboxRom_81;
  wire       [7:0]    sboxRom_82;
  wire       [7:0]    sboxRom_83;
  wire       [7:0]    sboxRom_84;
  wire       [7:0]    sboxRom_85;
  wire       [7:0]    sboxRom_86;
  wire       [7:0]    sboxRom_87;
  wire       [7:0]    sboxRom_88;
  wire       [7:0]    sboxRom_89;
  wire       [7:0]    sboxRom_90;
  wire       [7:0]    sboxRom_91;
  wire       [7:0]    sboxRom_92;
  wire       [7:0]    sboxRom_93;
  wire       [7:0]    sboxRom_94;
  wire       [7:0]    sboxRom_95;
  wire       [7:0]    sboxRom_96;
  wire       [7:0]    sboxRom_97;
  wire       [7:0]    sboxRom_98;
  wire       [7:0]    sboxRom_99;
  wire       [7:0]    sboxRom_100;
  wire       [7:0]    sboxRom_101;
  wire       [7:0]    sboxRom_102;
  wire       [7:0]    sboxRom_103;
  wire       [7:0]    sboxRom_104;
  wire       [7:0]    sboxRom_105;
  wire       [7:0]    sboxRom_106;
  wire       [7:0]    sboxRom_107;
  wire       [7:0]    sboxRom_108;
  wire       [7:0]    sboxRom_109;
  wire       [7:0]    sboxRom_110;
  wire       [7:0]    sboxRom_111;
  wire       [7:0]    sboxRom_112;
  wire       [7:0]    sboxRom_113;
  wire       [7:0]    sboxRom_114;
  wire       [7:0]    sboxRom_115;
  wire       [7:0]    sboxRom_116;
  wire       [7:0]    sboxRom_117;
  wire       [7:0]    sboxRom_118;
  wire       [7:0]    sboxRom_119;
  wire       [7:0]    sboxRom_120;
  wire       [7:0]    sboxRom_121;
  wire       [7:0]    sboxRom_122;
  wire       [7:0]    sboxRom_123;
  wire       [7:0]    sboxRom_124;
  wire       [7:0]    sboxRom_125;
  wire       [7:0]    sboxRom_126;
  wire       [7:0]    sboxRom_127;
  wire       [7:0]    sboxRom_128;
  wire       [7:0]    sboxRom_129;
  wire       [7:0]    sboxRom_130;
  wire       [7:0]    sboxRom_131;
  wire       [7:0]    sboxRom_132;
  wire       [7:0]    sboxRom_133;
  wire       [7:0]    sboxRom_134;
  wire       [7:0]    sboxRom_135;
  wire       [7:0]    sboxRom_136;
  wire       [7:0]    sboxRom_137;
  wire       [7:0]    sboxRom_138;
  wire       [7:0]    sboxRom_139;
  wire       [7:0]    sboxRom_140;
  wire       [7:0]    sboxRom_141;
  wire       [7:0]    sboxRom_142;
  wire       [7:0]    sboxRom_143;
  wire       [7:0]    sboxRom_144;
  wire       [7:0]    sboxRom_145;
  wire       [7:0]    sboxRom_146;
  wire       [7:0]    sboxRom_147;
  wire       [7:0]    sboxRom_148;
  wire       [7:0]    sboxRom_149;
  wire       [7:0]    sboxRom_150;
  wire       [7:0]    sboxRom_151;
  wire       [7:0]    sboxRom_152;
  wire       [7:0]    sboxRom_153;
  wire       [7:0]    sboxRom_154;
  wire       [7:0]    sboxRom_155;
  wire       [7:0]    sboxRom_156;
  wire       [7:0]    sboxRom_157;
  wire       [7:0]    sboxRom_158;
  wire       [7:0]    sboxRom_159;
  wire       [7:0]    sboxRom_160;
  wire       [7:0]    sboxRom_161;
  wire       [7:0]    sboxRom_162;
  wire       [7:0]    sboxRom_163;
  wire       [7:0]    sboxRom_164;
  wire       [7:0]    sboxRom_165;
  wire       [7:0]    sboxRom_166;
  wire       [7:0]    sboxRom_167;
  wire       [7:0]    sboxRom_168;
  wire       [7:0]    sboxRom_169;
  wire       [7:0]    sboxRom_170;
  wire       [7:0]    sboxRom_171;
  wire       [7:0]    sboxRom_172;
  wire       [7:0]    sboxRom_173;
  wire       [7:0]    sboxRom_174;
  wire       [7:0]    sboxRom_175;
  wire       [7:0]    sboxRom_176;
  wire       [7:0]    sboxRom_177;
  wire       [7:0]    sboxRom_178;
  wire       [7:0]    sboxRom_179;
  wire       [7:0]    sboxRom_180;
  wire       [7:0]    sboxRom_181;
  wire       [7:0]    sboxRom_182;
  wire       [7:0]    sboxRom_183;
  wire       [7:0]    sboxRom_184;
  wire       [7:0]    sboxRom_185;
  wire       [7:0]    sboxRom_186;
  wire       [7:0]    sboxRom_187;
  wire       [7:0]    sboxRom_188;
  wire       [7:0]    sboxRom_189;
  wire       [7:0]    sboxRom_190;
  wire       [7:0]    sboxRom_191;
  wire       [7:0]    sboxRom_192;
  wire       [7:0]    sboxRom_193;
  wire       [7:0]    sboxRom_194;
  wire       [7:0]    sboxRom_195;
  wire       [7:0]    sboxRom_196;
  wire       [7:0]    sboxRom_197;
  wire       [7:0]    sboxRom_198;
  wire       [7:0]    sboxRom_199;
  wire       [7:0]    sboxRom_200;
  wire       [7:0]    sboxRom_201;
  wire       [7:0]    sboxRom_202;
  wire       [7:0]    sboxRom_203;
  wire       [7:0]    sboxRom_204;
  wire       [7:0]    sboxRom_205;
  wire       [7:0]    sboxRom_206;
  wire       [7:0]    sboxRom_207;
  wire       [7:0]    sboxRom_208;
  wire       [7:0]    sboxRom_209;
  wire       [7:0]    sboxRom_210;
  wire       [7:0]    sboxRom_211;
  wire       [7:0]    sboxRom_212;
  wire       [7:0]    sboxRom_213;
  wire       [7:0]    sboxRom_214;
  wire       [7:0]    sboxRom_215;
  wire       [7:0]    sboxRom_216;
  wire       [7:0]    sboxRom_217;
  wire       [7:0]    sboxRom_218;
  wire       [7:0]    sboxRom_219;
  wire       [7:0]    sboxRom_220;
  wire       [7:0]    sboxRom_221;
  wire       [7:0]    sboxRom_222;
  wire       [7:0]    sboxRom_223;
  wire       [7:0]    sboxRom_224;
  wire       [7:0]    sboxRom_225;
  wire       [7:0]    sboxRom_226;
  wire       [7:0]    sboxRom_227;
  wire       [7:0]    sboxRom_228;
  wire       [7:0]    sboxRom_229;
  wire       [7:0]    sboxRom_230;
  wire       [7:0]    sboxRom_231;
  wire       [7:0]    sboxRom_232;
  wire       [7:0]    sboxRom_233;
  wire       [7:0]    sboxRom_234;
  wire       [7:0]    sboxRom_235;
  wire       [7:0]    sboxRom_236;
  wire       [7:0]    sboxRom_237;
  wire       [7:0]    sboxRom_238;
  wire       [7:0]    sboxRom_239;
  wire       [7:0]    sboxRom_240;
  wire       [7:0]    sboxRom_241;
  wire       [7:0]    sboxRom_242;
  wire       [7:0]    sboxRom_243;
  wire       [7:0]    sboxRom_244;
  wire       [7:0]    sboxRom_245;
  wire       [7:0]    sboxRom_246;
  wire       [7:0]    sboxRom_247;
  wire       [7:0]    sboxRom_248;
  wire       [7:0]    sboxRom_249;
  wire       [7:0]    sboxRom_250;
  wire       [7:0]    sboxRom_251;
  wire       [7:0]    sboxRom_252;
  wire       [7:0]    sboxRom_253;
  wire       [7:0]    sboxRom_254;
  wire       [7:0]    sboxRom_255;
  wire       [7:0]    rcon_0;
  wire       [7:0]    rcon_1;
  wire       [7:0]    rcon_2;
  wire       [7:0]    rcon_3;
  wire       [7:0]    rcon_4;
  wire       [7:0]    rcon_5;
  wire       [7:0]    rcon_6;
  wire       [7:0]    rcon_7;
  wire       [7:0]    rcon_8;
  wire       [7:0]    rcon_9;
  reg        [127:0]  stateReg;
  reg        [31:0]   roundKeyReg_0;
  reg        [31:0]   roundKeyReg_1;
  reg        [31:0]   roundKeyReg_2;
  reg        [31:0]   roundKeyReg_3;
  reg        [3:0]    roundCount;
  reg                 running;
  reg        [3:0]    rconCounter;
  reg        [127:0]  newStateComb;
  reg        [127:0]  rkBitsUsedComb;
  wire       [7:0]    invSboxRom_0;
  wire       [7:0]    invSboxRom_1;
  wire       [7:0]    invSboxRom_2;
  wire       [7:0]    invSboxRom_3;
  wire       [7:0]    invSboxRom_4;
  wire       [7:0]    invSboxRom_5;
  wire       [7:0]    invSboxRom_6;
  wire       [7:0]    invSboxRom_7;
  wire       [7:0]    invSboxRom_8;
  wire       [7:0]    invSboxRom_9;
  wire       [7:0]    invSboxRom_10;
  wire       [7:0]    invSboxRom_11;
  wire       [7:0]    invSboxRom_12;
  wire       [7:0]    invSboxRom_13;
  wire       [7:0]    invSboxRom_14;
  wire       [7:0]    invSboxRom_15;
  wire       [7:0]    invSboxRom_16;
  wire       [7:0]    invSboxRom_17;
  wire       [7:0]    invSboxRom_18;
  wire       [7:0]    invSboxRom_19;
  wire       [7:0]    invSboxRom_20;
  wire       [7:0]    invSboxRom_21;
  wire       [7:0]    invSboxRom_22;
  wire       [7:0]    invSboxRom_23;
  wire       [7:0]    invSboxRom_24;
  wire       [7:0]    invSboxRom_25;
  wire       [7:0]    invSboxRom_26;
  wire       [7:0]    invSboxRom_27;
  wire       [7:0]    invSboxRom_28;
  wire       [7:0]    invSboxRom_29;
  wire       [7:0]    invSboxRom_30;
  wire       [7:0]    invSboxRom_31;
  wire       [7:0]    invSboxRom_32;
  wire       [7:0]    invSboxRom_33;
  wire       [7:0]    invSboxRom_34;
  wire       [7:0]    invSboxRom_35;
  wire       [7:0]    invSboxRom_36;
  wire       [7:0]    invSboxRom_37;
  wire       [7:0]    invSboxRom_38;
  wire       [7:0]    invSboxRom_39;
  wire       [7:0]    invSboxRom_40;
  wire       [7:0]    invSboxRom_41;
  wire       [7:0]    invSboxRom_42;
  wire       [7:0]    invSboxRom_43;
  wire       [7:0]    invSboxRom_44;
  wire       [7:0]    invSboxRom_45;
  wire       [7:0]    invSboxRom_46;
  wire       [7:0]    invSboxRom_47;
  wire       [7:0]    invSboxRom_48;
  wire       [7:0]    invSboxRom_49;
  wire       [7:0]    invSboxRom_50;
  wire       [7:0]    invSboxRom_51;
  wire       [7:0]    invSboxRom_52;
  wire       [7:0]    invSboxRom_53;
  wire       [7:0]    invSboxRom_54;
  wire       [7:0]    invSboxRom_55;
  wire       [7:0]    invSboxRom_56;
  wire       [7:0]    invSboxRom_57;
  wire       [7:0]    invSboxRom_58;
  wire       [7:0]    invSboxRom_59;
  wire       [7:0]    invSboxRom_60;
  wire       [7:0]    invSboxRom_61;
  wire       [7:0]    invSboxRom_62;
  wire       [7:0]    invSboxRom_63;
  wire       [7:0]    invSboxRom_64;
  wire       [7:0]    invSboxRom_65;
  wire       [7:0]    invSboxRom_66;
  wire       [7:0]    invSboxRom_67;
  wire       [7:0]    invSboxRom_68;
  wire       [7:0]    invSboxRom_69;
  wire       [7:0]    invSboxRom_70;
  wire       [7:0]    invSboxRom_71;
  wire       [7:0]    invSboxRom_72;
  wire       [7:0]    invSboxRom_73;
  wire       [7:0]    invSboxRom_74;
  wire       [7:0]    invSboxRom_75;
  wire       [7:0]    invSboxRom_76;
  wire       [7:0]    invSboxRom_77;
  wire       [7:0]    invSboxRom_78;
  wire       [7:0]    invSboxRom_79;
  wire       [7:0]    invSboxRom_80;
  wire       [7:0]    invSboxRom_81;
  wire       [7:0]    invSboxRom_82;
  wire       [7:0]    invSboxRom_83;
  wire       [7:0]    invSboxRom_84;
  wire       [7:0]    invSboxRom_85;
  wire       [7:0]    invSboxRom_86;
  wire       [7:0]    invSboxRom_87;
  wire       [7:0]    invSboxRom_88;
  wire       [7:0]    invSboxRom_89;
  wire       [7:0]    invSboxRom_90;
  wire       [7:0]    invSboxRom_91;
  wire       [7:0]    invSboxRom_92;
  wire       [7:0]    invSboxRom_93;
  wire       [7:0]    invSboxRom_94;
  wire       [7:0]    invSboxRom_95;
  wire       [7:0]    invSboxRom_96;
  wire       [7:0]    invSboxRom_97;
  wire       [7:0]    invSboxRom_98;
  wire       [7:0]    invSboxRom_99;
  wire       [7:0]    invSboxRom_100;
  wire       [7:0]    invSboxRom_101;
  wire       [7:0]    invSboxRom_102;
  wire       [7:0]    invSboxRom_103;
  wire       [7:0]    invSboxRom_104;
  wire       [7:0]    invSboxRom_105;
  wire       [7:0]    invSboxRom_106;
  wire       [7:0]    invSboxRom_107;
  wire       [7:0]    invSboxRom_108;
  wire       [7:0]    invSboxRom_109;
  wire       [7:0]    invSboxRom_110;
  wire       [7:0]    invSboxRom_111;
  wire       [7:0]    invSboxRom_112;
  wire       [7:0]    invSboxRom_113;
  wire       [7:0]    invSboxRom_114;
  wire       [7:0]    invSboxRom_115;
  wire       [7:0]    invSboxRom_116;
  wire       [7:0]    invSboxRom_117;
  wire       [7:0]    invSboxRom_118;
  wire       [7:0]    invSboxRom_119;
  wire       [7:0]    invSboxRom_120;
  wire       [7:0]    invSboxRom_121;
  wire       [7:0]    invSboxRom_122;
  wire       [7:0]    invSboxRom_123;
  wire       [7:0]    invSboxRom_124;
  wire       [7:0]    invSboxRom_125;
  wire       [7:0]    invSboxRom_126;
  wire       [7:0]    invSboxRom_127;
  wire       [7:0]    invSboxRom_128;
  wire       [7:0]    invSboxRom_129;
  wire       [7:0]    invSboxRom_130;
  wire       [7:0]    invSboxRom_131;
  wire       [7:0]    invSboxRom_132;
  wire       [7:0]    invSboxRom_133;
  wire       [7:0]    invSboxRom_134;
  wire       [7:0]    invSboxRom_135;
  wire       [7:0]    invSboxRom_136;
  wire       [7:0]    invSboxRom_137;
  wire       [7:0]    invSboxRom_138;
  wire       [7:0]    invSboxRom_139;
  wire       [7:0]    invSboxRom_140;
  wire       [7:0]    invSboxRom_141;
  wire       [7:0]    invSboxRom_142;
  wire       [7:0]    invSboxRom_143;
  wire       [7:0]    invSboxRom_144;
  wire       [7:0]    invSboxRom_145;
  wire       [7:0]    invSboxRom_146;
  wire       [7:0]    invSboxRom_147;
  wire       [7:0]    invSboxRom_148;
  wire       [7:0]    invSboxRom_149;
  wire       [7:0]    invSboxRom_150;
  wire       [7:0]    invSboxRom_151;
  wire       [7:0]    invSboxRom_152;
  wire       [7:0]    invSboxRom_153;
  wire       [7:0]    invSboxRom_154;
  wire       [7:0]    invSboxRom_155;
  wire       [7:0]    invSboxRom_156;
  wire       [7:0]    invSboxRom_157;
  wire       [7:0]    invSboxRom_158;
  wire       [7:0]    invSboxRom_159;
  wire       [7:0]    invSboxRom_160;
  wire       [7:0]    invSboxRom_161;
  wire       [7:0]    invSboxRom_162;
  wire       [7:0]    invSboxRom_163;
  wire       [7:0]    invSboxRom_164;
  wire       [7:0]    invSboxRom_165;
  wire       [7:0]    invSboxRom_166;
  wire       [7:0]    invSboxRom_167;
  wire       [7:0]    invSboxRom_168;
  wire       [7:0]    invSboxRom_169;
  wire       [7:0]    invSboxRom_170;
  wire       [7:0]    invSboxRom_171;
  wire       [7:0]    invSboxRom_172;
  wire       [7:0]    invSboxRom_173;
  wire       [7:0]    invSboxRom_174;
  wire       [7:0]    invSboxRom_175;
  wire       [7:0]    invSboxRom_176;
  wire       [7:0]    invSboxRom_177;
  wire       [7:0]    invSboxRom_178;
  wire       [7:0]    invSboxRom_179;
  wire       [7:0]    invSboxRom_180;
  wire       [7:0]    invSboxRom_181;
  wire       [7:0]    invSboxRom_182;
  wire       [7:0]    invSboxRom_183;
  wire       [7:0]    invSboxRom_184;
  wire       [7:0]    invSboxRom_185;
  wire       [7:0]    invSboxRom_186;
  wire       [7:0]    invSboxRom_187;
  wire       [7:0]    invSboxRom_188;
  wire       [7:0]    invSboxRom_189;
  wire       [7:0]    invSboxRom_190;
  wire       [7:0]    invSboxRom_191;
  wire       [7:0]    invSboxRom_192;
  wire       [7:0]    invSboxRom_193;
  wire       [7:0]    invSboxRom_194;
  wire       [7:0]    invSboxRom_195;
  wire       [7:0]    invSboxRom_196;
  wire       [7:0]    invSboxRom_197;
  wire       [7:0]    invSboxRom_198;
  wire       [7:0]    invSboxRom_199;
  wire       [7:0]    invSboxRom_200;
  wire       [7:0]    invSboxRom_201;
  wire       [7:0]    invSboxRom_202;
  wire       [7:0]    invSboxRom_203;
  wire       [7:0]    invSboxRom_204;
  wire       [7:0]    invSboxRom_205;
  wire       [7:0]    invSboxRom_206;
  wire       [7:0]    invSboxRom_207;
  wire       [7:0]    invSboxRom_208;
  wire       [7:0]    invSboxRom_209;
  wire       [7:0]    invSboxRom_210;
  wire       [7:0]    invSboxRom_211;
  wire       [7:0]    invSboxRom_212;
  wire       [7:0]    invSboxRom_213;
  wire       [7:0]    invSboxRom_214;
  wire       [7:0]    invSboxRom_215;
  wire       [7:0]    invSboxRom_216;
  wire       [7:0]    invSboxRom_217;
  wire       [7:0]    invSboxRom_218;
  wire       [7:0]    invSboxRom_219;
  wire       [7:0]    invSboxRom_220;
  wire       [7:0]    invSboxRom_221;
  wire       [7:0]    invSboxRom_222;
  wire       [7:0]    invSboxRom_223;
  wire       [7:0]    invSboxRom_224;
  wire       [7:0]    invSboxRom_225;
  wire       [7:0]    invSboxRom_226;
  wire       [7:0]    invSboxRom_227;
  wire       [7:0]    invSboxRom_228;
  wire       [7:0]    invSboxRom_229;
  wire       [7:0]    invSboxRom_230;
  wire       [7:0]    invSboxRom_231;
  wire       [7:0]    invSboxRom_232;
  wire       [7:0]    invSboxRom_233;
  wire       [7:0]    invSboxRom_234;
  wire       [7:0]    invSboxRom_235;
  wire       [7:0]    invSboxRom_236;
  wire       [7:0]    invSboxRom_237;
  wire       [7:0]    invSboxRom_238;
  wire       [7:0]    invSboxRom_239;
  wire       [7:0]    invSboxRom_240;
  wire       [7:0]    invSboxRom_241;
  wire       [7:0]    invSboxRom_242;
  wire       [7:0]    invSboxRom_243;
  wire       [7:0]    invSboxRom_244;
  wire       [7:0]    invSboxRom_245;
  wire       [7:0]    invSboxRom_246;
  wire       [7:0]    invSboxRom_247;
  wire       [7:0]    invSboxRom_248;
  wire       [7:0]    invSboxRom_249;
  wire       [7:0]    invSboxRom_250;
  wire       [7:0]    invSboxRom_251;
  wire       [7:0]    invSboxRom_252;
  wire       [7:0]    invSboxRom_253;
  wire       [7:0]    invSboxRom_254;
  wire       [7:0]    invSboxRom_255;
  reg                 precomputeRunning;
  reg        [3:0]    precomputeCounter;
  reg        [31:0]   initKeyWords_0;
  reg        [31:0]   initKeyWords_1;
  reg        [31:0]   initKeyWords_2;
  reg        [31:0]   initKeyWords_3;
  reg        [7:0]    invShifted_0;
  reg        [7:0]    invShifted_1;
  reg        [7:0]    invShifted_2;
  reg        [7:0]    invShifted_3;
  reg        [7:0]    invShifted_4;
  reg        [7:0]    invShifted_5;
  reg        [7:0]    invShifted_6;
  reg        [7:0]    invShifted_7;
  reg        [7:0]    invShifted_8;
  reg        [7:0]    invShifted_9;
  reg        [7:0]    invShifted_10;
  reg        [7:0]    invShifted_11;
  reg        [7:0]    invShifted_12;
  reg        [7:0]    invShifted_13;
  reg        [7:0]    invShifted_14;
  reg        [7:0]    invShifted_15;
  reg        [7:0]    invSub_0;
  reg        [7:0]    invSub_1;
  reg        [7:0]    invSub_2;
  reg        [7:0]    invSub_3;
  reg        [7:0]    invSub_4;
  reg        [7:0]    invSub_5;
  reg        [7:0]    invSub_6;
  reg        [7:0]    invSub_7;
  reg        [7:0]    invSub_8;
  reg        [7:0]    invSub_9;
  reg        [7:0]    invSub_10;
  reg        [7:0]    invSub_11;
  reg        [7:0]    invSub_12;
  reg        [7:0]    invSub_13;
  reg        [7:0]    invSub_14;
  reg        [7:0]    invSub_15;
  reg        [7:0]    invMixed_0;
  reg        [7:0]    invMixed_1;
  reg        [7:0]    invMixed_2;
  reg        [7:0]    invMixed_3;
  reg        [7:0]    invMixed_4;
  reg        [7:0]    invMixed_5;
  reg        [7:0]    invMixed_6;
  reg        [7:0]    invMixed_7;
  reg        [7:0]    invMixed_8;
  reg        [7:0]    invMixed_9;
  reg        [7:0]    invMixed_10;
  reg        [7:0]    invMixed_11;
  reg        [7:0]    invMixed_12;
  reg        [7:0]    invMixed_13;
  reg        [7:0]    invMixed_14;
  reg        [7:0]    invMixed_15;
  wire                when_AES128_l230;
  wire       [31:0]   _zz_stateReg;
  wire       [31:0]   _zz_stateReg_1;
  wire       [31:0]   _zz_stateReg_2;
  wire       [31:0]   _zz_stateReg_3;
  wire       [7:0]    _zz_stateReg_4;
  wire       [7:0]    _zz_stateReg_5;
  wire       [7:0]    _zz_stateReg_6;
  wire       [7:0]    _zz_stateReg_7;
  wire       [7:0]    _zz_stateReg_8;
  wire       [7:0]    _zz_stateReg_9;
  wire       [7:0]    _zz_stateReg_10;
  wire       [7:0]    _zz_stateReg_11;
  wire       [7:0]    _zz_stateReg_12;
  wire       [7:0]    _zz_stateReg_13;
  wire       [7:0]    _zz_stateReg_14;
  wire       [7:0]    _zz_stateReg_15;
  wire       [7:0]    _zz_stateReg_16;
  wire       [7:0]    _zz_stateReg_17;
  wire       [7:0]    _zz_stateReg_18;
  wire       [7:0]    _zz_stateReg_19;
  reg        [7:0]    _zz_stateReg_20;
  reg        [7:0]    _zz_stateReg_21;
  reg        [7:0]    _zz_stateReg_22;
  reg        [7:0]    _zz_stateReg_23;
  reg        [7:0]    _zz_stateReg_24;
  reg        [7:0]    _zz_stateReg_25;
  reg        [7:0]    _zz_stateReg_26;
  reg        [7:0]    _zz_stateReg_27;
  reg        [7:0]    _zz_stateReg_28;
  reg        [7:0]    _zz_stateReg_29;
  reg        [7:0]    _zz_stateReg_30;
  reg        [7:0]    _zz_stateReg_31;
  reg        [7:0]    _zz_stateReg_32;
  reg        [7:0]    _zz_stateReg_33;
  reg        [7:0]    _zz_stateReg_34;
  reg        [7:0]    _zz_stateReg_35;
  wire                when_AES128_l272;
  wire       [7:0]    _zz_stateReg_36;
  wire       [7:0]    _zz_stateReg_37;
  wire       [7:0]    _zz_stateReg_38;
  wire       [7:0]    _zz_stateReg_39;
  wire       [7:0]    _zz_stateReg_40;
  wire       [7:0]    _zz_stateReg_41;
  wire       [7:0]    _zz_stateReg_42;
  wire       [7:0]    _zz_stateReg_43;
  wire       [7:0]    _zz_stateReg_44;
  wire       [7:0]    _zz_stateReg_45;
  wire       [7:0]    _zz_stateReg_46;
  wire       [7:0]    _zz_stateReg_47;
  wire       [7:0]    _zz_stateReg_48;
  wire       [7:0]    _zz_stateReg_49;
  wire       [7:0]    _zz_stateReg_50;
  wire       [7:0]    _zz_stateReg_51;
  wire       [7:0]    _zz_stateReg_52;
  wire       [7:0]    _zz_stateReg_53;
  wire       [7:0]    _zz_stateReg_54;
  wire       [7:0]    _zz_stateReg_55;
  wire       [7:0]    _zz_stateReg_56;
  wire       [7:0]    _zz_stateReg_57;
  wire       [7:0]    _zz_stateReg_58;
  wire       [7:0]    _zz_stateReg_59;
  wire       [7:0]    _zz_stateReg_60;
  wire       [7:0]    _zz_stateReg_61;
  wire       [7:0]    _zz_stateReg_62;
  wire       [7:0]    _zz_stateReg_63;
  wire       [7:0]    _zz_stateReg_64;
  wire       [7:0]    _zz_stateReg_65;
  wire       [7:0]    _zz_stateReg_66;
  wire       [7:0]    _zz_stateReg_67;
  wire       [127:0]  _zz_stateReg_68;
  wire       [7:0]    _zz_roundKeyReg_0;
  wire       [31:0]   _zz_roundKeyReg_0_1;
  wire       [31:0]   _zz_roundKeyReg_0_2;
  wire       [31:0]   _zz_roundKeyReg_1;
  wire       [31:0]   _zz_roundKeyReg_2;
  wire       [31:0]   _zz_roundKeyReg_3;
  wire       [127:0]  _zz_stateReg_69;
  wire                when_AES128_l307;
  wire                when_AES128_l313;
  wire       [31:0]   _zz_roundKeyReg_0_3;
  wire       [31:0]   _zz_roundKeyReg_1_1;
  wire       [31:0]   _zz_roundKeyReg_2_1;
  wire       [31:0]   _zz_roundKeyReg_3_1;
  wire       [31:0]   _zz_stateReg_70;
  wire       [31:0]   _zz_stateReg_71;
  wire       [31:0]   _zz_stateReg_72;
  wire       [31:0]   _zz_stateReg_73;
  wire       [31:0]   _zz_stateReg_74;
  wire                when_AES128_l328;
  wire       [31:0]   _zz_roundKeyReg_3_2;
  wire       [31:0]   _zz_roundKeyReg_2_2;
  wire       [31:0]   _zz_roundKeyReg_1_2;
  wire       [31:0]   _zz_roundKeyReg_0_4;
  wire       [31:0]   _zz_roundKeyReg_0_5;
  wire       [127:0]  _zz_invMixed_0;
  wire       [7:0]    _zz_invMixed_0_1;
  wire       [7:0]    _zz_invMixed_0_2;
  wire       [7:0]    _zz_invMixed_0_3;
  wire       [7:0]    _zz_invMixed_0_4;
  wire       [7:0]    _zz_invMixed_4;
  wire       [7:0]    _zz_invMixed_4_1;
  wire       [7:0]    _zz_invMixed_4_2;
  wire       [7:0]    _zz_invMixed_4_3;
  wire       [7:0]    _zz_invMixed_8;
  wire       [7:0]    _zz_invMixed_8_1;
  wire       [7:0]    _zz_invMixed_8_2;
  wire       [7:0]    _zz_invMixed_8_3;
  wire       [7:0]    _zz_invMixed_12;
  wire       [7:0]    _zz_invMixed_12_1;
  wire       [7:0]    _zz_invMixed_12_2;
  wire       [7:0]    _zz_invMixed_12_3;
  wire                when_AES128_l370;
  wire       [7:0]    _zz_invMixed_0_5;
  wire       [7:0]    _zz_invMixed_0_6;
  wire       [7:0]    _zz_invMixed_0_7;
  wire       [7:0]    _zz_invMixed_0_8;
  wire       [7:0]    _zz_invMixed_0_9;
  wire       [7:0]    _zz_invMixed_0_10;
  wire       [7:0]    _zz_invMixed_0_11;
  wire       [7:0]    _zz_invMixed_0_12;
  wire       [7:0]    _zz_invMixed_0_13;
  wire       [7:0]    _zz_invMixed_0_14;
  wire       [7:0]    _zz_invMixed_0_15;
  wire       [7:0]    _zz_invMixed_0_16;
  wire       [7:0]    _zz_invMixed_0_17;
  wire       [7:0]    _zz_invMixed_0_18;
  wire       [7:0]    _zz_invMixed_0_19;
  wire       [7:0]    _zz_invMixed_0_20;
  wire       [7:0]    _zz_invMixed_0_21;
  wire       [7:0]    _zz_invMixed_0_22;
  wire       [7:0]    _zz_invMixed_0_23;
  wire       [7:0]    _zz_invMixed_0_24;
  wire       [7:0]    _zz_invMixed_0_25;
  wire       [7:0]    _zz_invMixed_0_26;
  wire       [7:0]    _zz_invMixed_0_27;
  wire       [7:0]    _zz_invMixed_0_28;
  wire       [7:0]    _zz_invMixed_0_29;
  wire       [7:0]    _zz_invMixed_0_30;
  wire       [7:0]    _zz_invMixed_0_31;
  wire       [7:0]    _zz_invMixed_0_32;
  wire       [7:0]    _zz_invMixed_1;
  wire       [7:0]    _zz_invMixed_1_1;
  wire       [7:0]    _zz_invMixed_1_2;
  wire       [7:0]    _zz_invMixed_1_3;
  wire       [7:0]    _zz_invMixed_1_4;
  wire       [7:0]    _zz_invMixed_1_5;
  wire       [7:0]    _zz_invMixed_1_6;
  wire       [7:0]    _zz_invMixed_1_7;
  wire       [7:0]    _zz_invMixed_1_8;
  wire       [7:0]    _zz_invMixed_1_9;
  wire       [7:0]    _zz_invMixed_1_10;
  wire       [7:0]    _zz_invMixed_1_11;
  wire       [7:0]    _zz_invMixed_1_12;
  wire       [7:0]    _zz_invMixed_1_13;
  wire       [7:0]    _zz_invMixed_1_14;
  wire       [7:0]    _zz_invMixed_1_15;
  wire       [7:0]    _zz_invMixed_1_16;
  wire       [7:0]    _zz_invMixed_1_17;
  wire       [7:0]    _zz_invMixed_1_18;
  wire       [7:0]    _zz_invMixed_1_19;
  wire       [7:0]    _zz_invMixed_1_20;
  wire       [7:0]    _zz_invMixed_1_21;
  wire       [7:0]    _zz_invMixed_1_22;
  wire       [7:0]    _zz_invMixed_1_23;
  wire       [7:0]    _zz_invMixed_1_24;
  wire       [7:0]    _zz_invMixed_1_25;
  wire       [7:0]    _zz_invMixed_1_26;
  wire       [7:0]    _zz_invMixed_1_27;
  wire       [7:0]    _zz_invMixed_2;
  wire       [7:0]    _zz_invMixed_2_1;
  wire       [7:0]    _zz_invMixed_2_2;
  wire       [7:0]    _zz_invMixed_2_3;
  wire       [7:0]    _zz_invMixed_2_4;
  wire       [7:0]    _zz_invMixed_2_5;
  wire       [7:0]    _zz_invMixed_2_6;
  wire       [7:0]    _zz_invMixed_2_7;
  wire       [7:0]    _zz_invMixed_2_8;
  wire       [7:0]    _zz_invMixed_2_9;
  wire       [7:0]    _zz_invMixed_2_10;
  wire       [7:0]    _zz_invMixed_2_11;
  wire       [7:0]    _zz_invMixed_2_12;
  wire       [7:0]    _zz_invMixed_2_13;
  wire       [7:0]    _zz_invMixed_2_14;
  wire       [7:0]    _zz_invMixed_2_15;
  wire       [7:0]    _zz_invMixed_2_16;
  wire       [7:0]    _zz_invMixed_2_17;
  wire       [7:0]    _zz_invMixed_2_18;
  wire       [7:0]    _zz_invMixed_2_19;
  wire       [7:0]    _zz_invMixed_2_20;
  wire       [7:0]    _zz_invMixed_2_21;
  wire       [7:0]    _zz_invMixed_2_22;
  wire       [7:0]    _zz_invMixed_2_23;
  wire       [7:0]    _zz_invMixed_2_24;
  wire       [7:0]    _zz_invMixed_2_25;
  wire       [7:0]    _zz_invMixed_2_26;
  wire       [7:0]    _zz_invMixed_2_27;
  wire       [7:0]    _zz_invMixed_3;
  wire       [7:0]    _zz_invMixed_3_1;
  wire       [7:0]    _zz_invMixed_3_2;
  wire       [7:0]    _zz_invMixed_3_3;
  wire       [7:0]    _zz_invMixed_3_4;
  wire       [7:0]    _zz_invMixed_3_5;
  wire       [7:0]    _zz_invMixed_3_6;
  wire       [7:0]    _zz_invMixed_3_7;
  wire       [7:0]    _zz_invMixed_3_8;
  wire       [7:0]    _zz_invMixed_3_9;
  wire       [7:0]    _zz_invMixed_3_10;
  wire       [7:0]    _zz_invMixed_3_11;
  wire       [7:0]    _zz_invMixed_3_12;
  wire       [7:0]    _zz_invMixed_3_13;
  wire       [7:0]    _zz_invMixed_3_14;
  wire       [7:0]    _zz_invMixed_3_15;
  wire       [7:0]    _zz_invMixed_3_16;
  wire       [7:0]    _zz_invMixed_3_17;
  wire       [7:0]    _zz_invMixed_3_18;
  wire       [7:0]    _zz_invMixed_3_19;
  wire       [7:0]    _zz_invMixed_3_20;
  wire       [7:0]    _zz_invMixed_3_21;
  wire       [7:0]    _zz_invMixed_3_22;
  wire       [7:0]    _zz_invMixed_3_23;
  wire       [7:0]    _zz_invMixed_3_24;
  wire       [7:0]    _zz_invMixed_3_25;
  wire       [7:0]    _zz_invMixed_3_26;
  wire       [7:0]    _zz_invMixed_3_27;
  wire       [7:0]    _zz_invMixed_4_4;
  wire       [7:0]    _zz_invMixed_4_5;
  wire       [7:0]    _zz_invMixed_4_6;
  wire       [7:0]    _zz_invMixed_4_7;
  wire       [7:0]    _zz_invMixed_4_8;
  wire       [7:0]    _zz_invMixed_4_9;
  wire       [7:0]    _zz_invMixed_4_10;
  wire       [7:0]    _zz_invMixed_4_11;
  wire       [7:0]    _zz_invMixed_4_12;
  wire       [7:0]    _zz_invMixed_4_13;
  wire       [7:0]    _zz_invMixed_4_14;
  wire       [7:0]    _zz_invMixed_4_15;
  wire       [7:0]    _zz_invMixed_4_16;
  wire       [7:0]    _zz_invMixed_4_17;
  wire       [7:0]    _zz_invMixed_4_18;
  wire       [7:0]    _zz_invMixed_4_19;
  wire       [7:0]    _zz_invMixed_4_20;
  wire       [7:0]    _zz_invMixed_4_21;
  wire       [7:0]    _zz_invMixed_4_22;
  wire       [7:0]    _zz_invMixed_4_23;
  wire       [7:0]    _zz_invMixed_4_24;
  wire       [7:0]    _zz_invMixed_4_25;
  wire       [7:0]    _zz_invMixed_4_26;
  wire       [7:0]    _zz_invMixed_4_27;
  wire       [7:0]    _zz_invMixed_4_28;
  wire       [7:0]    _zz_invMixed_4_29;
  wire       [7:0]    _zz_invMixed_4_30;
  wire       [7:0]    _zz_invMixed_4_31;
  wire       [7:0]    _zz_invMixed_5;
  wire       [7:0]    _zz_invMixed_5_1;
  wire       [7:0]    _zz_invMixed_5_2;
  wire       [7:0]    _zz_invMixed_5_3;
  wire       [7:0]    _zz_invMixed_5_4;
  wire       [7:0]    _zz_invMixed_5_5;
  wire       [7:0]    _zz_invMixed_5_6;
  wire       [7:0]    _zz_invMixed_5_7;
  wire       [7:0]    _zz_invMixed_5_8;
  wire       [7:0]    _zz_invMixed_5_9;
  wire       [7:0]    _zz_invMixed_5_10;
  wire       [7:0]    _zz_invMixed_5_11;
  wire       [7:0]    _zz_invMixed_5_12;
  wire       [7:0]    _zz_invMixed_5_13;
  wire       [7:0]    _zz_invMixed_5_14;
  wire       [7:0]    _zz_invMixed_5_15;
  wire       [7:0]    _zz_invMixed_5_16;
  wire       [7:0]    _zz_invMixed_5_17;
  wire       [7:0]    _zz_invMixed_5_18;
  wire       [7:0]    _zz_invMixed_5_19;
  wire       [7:0]    _zz_invMixed_5_20;
  wire       [7:0]    _zz_invMixed_5_21;
  wire       [7:0]    _zz_invMixed_5_22;
  wire       [7:0]    _zz_invMixed_5_23;
  wire       [7:0]    _zz_invMixed_5_24;
  wire       [7:0]    _zz_invMixed_5_25;
  wire       [7:0]    _zz_invMixed_5_26;
  wire       [7:0]    _zz_invMixed_5_27;
  wire       [7:0]    _zz_invMixed_6;
  wire       [7:0]    _zz_invMixed_6_1;
  wire       [7:0]    _zz_invMixed_6_2;
  wire       [7:0]    _zz_invMixed_6_3;
  wire       [7:0]    _zz_invMixed_6_4;
  wire       [7:0]    _zz_invMixed_6_5;
  wire       [7:0]    _zz_invMixed_6_6;
  wire       [7:0]    _zz_invMixed_6_7;
  wire       [7:0]    _zz_invMixed_6_8;
  wire       [7:0]    _zz_invMixed_6_9;
  wire       [7:0]    _zz_invMixed_6_10;
  wire       [7:0]    _zz_invMixed_6_11;
  wire       [7:0]    _zz_invMixed_6_12;
  wire       [7:0]    _zz_invMixed_6_13;
  wire       [7:0]    _zz_invMixed_6_14;
  wire       [7:0]    _zz_invMixed_6_15;
  wire       [7:0]    _zz_invMixed_6_16;
  wire       [7:0]    _zz_invMixed_6_17;
  wire       [7:0]    _zz_invMixed_6_18;
  wire       [7:0]    _zz_invMixed_6_19;
  wire       [7:0]    _zz_invMixed_6_20;
  wire       [7:0]    _zz_invMixed_6_21;
  wire       [7:0]    _zz_invMixed_6_22;
  wire       [7:0]    _zz_invMixed_6_23;
  wire       [7:0]    _zz_invMixed_6_24;
  wire       [7:0]    _zz_invMixed_6_25;
  wire       [7:0]    _zz_invMixed_6_26;
  wire       [7:0]    _zz_invMixed_6_27;
  wire       [7:0]    _zz_invMixed_7;
  wire       [7:0]    _zz_invMixed_7_1;
  wire       [7:0]    _zz_invMixed_7_2;
  wire       [7:0]    _zz_invMixed_7_3;
  wire       [7:0]    _zz_invMixed_7_4;
  wire       [7:0]    _zz_invMixed_7_5;
  wire       [7:0]    _zz_invMixed_7_6;
  wire       [7:0]    _zz_invMixed_7_7;
  wire       [7:0]    _zz_invMixed_7_8;
  wire       [7:0]    _zz_invMixed_7_9;
  wire       [7:0]    _zz_invMixed_7_10;
  wire       [7:0]    _zz_invMixed_7_11;
  wire       [7:0]    _zz_invMixed_7_12;
  wire       [7:0]    _zz_invMixed_7_13;
  wire       [7:0]    _zz_invMixed_7_14;
  wire       [7:0]    _zz_invMixed_7_15;
  wire       [7:0]    _zz_invMixed_7_16;
  wire       [7:0]    _zz_invMixed_7_17;
  wire       [7:0]    _zz_invMixed_7_18;
  wire       [7:0]    _zz_invMixed_7_19;
  wire       [7:0]    _zz_invMixed_7_20;
  wire       [7:0]    _zz_invMixed_7_21;
  wire       [7:0]    _zz_invMixed_7_22;
  wire       [7:0]    _zz_invMixed_7_23;
  wire       [7:0]    _zz_invMixed_7_24;
  wire       [7:0]    _zz_invMixed_7_25;
  wire       [7:0]    _zz_invMixed_7_26;
  wire       [7:0]    _zz_invMixed_7_27;
  wire       [7:0]    _zz_invMixed_8_4;
  wire       [7:0]    _zz_invMixed_8_5;
  wire       [7:0]    _zz_invMixed_8_6;
  wire       [7:0]    _zz_invMixed_8_7;
  wire       [7:0]    _zz_invMixed_8_8;
  wire       [7:0]    _zz_invMixed_8_9;
  wire       [7:0]    _zz_invMixed_8_10;
  wire       [7:0]    _zz_invMixed_8_11;
  wire       [7:0]    _zz_invMixed_8_12;
  wire       [7:0]    _zz_invMixed_8_13;
  wire       [7:0]    _zz_invMixed_8_14;
  wire       [7:0]    _zz_invMixed_8_15;
  wire       [7:0]    _zz_invMixed_8_16;
  wire       [7:0]    _zz_invMixed_8_17;
  wire       [7:0]    _zz_invMixed_8_18;
  wire       [7:0]    _zz_invMixed_8_19;
  wire       [7:0]    _zz_invMixed_8_20;
  wire       [7:0]    _zz_invMixed_8_21;
  wire       [7:0]    _zz_invMixed_8_22;
  wire       [7:0]    _zz_invMixed_8_23;
  wire       [7:0]    _zz_invMixed_8_24;
  wire       [7:0]    _zz_invMixed_8_25;
  wire       [7:0]    _zz_invMixed_8_26;
  wire       [7:0]    _zz_invMixed_8_27;
  wire       [7:0]    _zz_invMixed_8_28;
  wire       [7:0]    _zz_invMixed_8_29;
  wire       [7:0]    _zz_invMixed_8_30;
  wire       [7:0]    _zz_invMixed_8_31;
  wire       [7:0]    _zz_invMixed_9;
  wire       [7:0]    _zz_invMixed_9_1;
  wire       [7:0]    _zz_invMixed_9_2;
  wire       [7:0]    _zz_invMixed_9_3;
  wire       [7:0]    _zz_invMixed_9_4;
  wire       [7:0]    _zz_invMixed_9_5;
  wire       [7:0]    _zz_invMixed_9_6;
  wire       [7:0]    _zz_invMixed_9_7;
  wire       [7:0]    _zz_invMixed_9_8;
  wire       [7:0]    _zz_invMixed_9_9;
  wire       [7:0]    _zz_invMixed_9_10;
  wire       [7:0]    _zz_invMixed_9_11;
  wire       [7:0]    _zz_invMixed_9_12;
  wire       [7:0]    _zz_invMixed_9_13;
  wire       [7:0]    _zz_invMixed_9_14;
  wire       [7:0]    _zz_invMixed_9_15;
  wire       [7:0]    _zz_invMixed_9_16;
  wire       [7:0]    _zz_invMixed_9_17;
  wire       [7:0]    _zz_invMixed_9_18;
  wire       [7:0]    _zz_invMixed_9_19;
  wire       [7:0]    _zz_invMixed_9_20;
  wire       [7:0]    _zz_invMixed_9_21;
  wire       [7:0]    _zz_invMixed_9_22;
  wire       [7:0]    _zz_invMixed_9_23;
  wire       [7:0]    _zz_invMixed_9_24;
  wire       [7:0]    _zz_invMixed_9_25;
  wire       [7:0]    _zz_invMixed_9_26;
  wire       [7:0]    _zz_invMixed_9_27;
  wire       [7:0]    _zz_invMixed_10;
  wire       [7:0]    _zz_invMixed_10_1;
  wire       [7:0]    _zz_invMixed_10_2;
  wire       [7:0]    _zz_invMixed_10_3;
  wire       [7:0]    _zz_invMixed_10_4;
  wire       [7:0]    _zz_invMixed_10_5;
  wire       [7:0]    _zz_invMixed_10_6;
  wire       [7:0]    _zz_invMixed_10_7;
  wire       [7:0]    _zz_invMixed_10_8;
  wire       [7:0]    _zz_invMixed_10_9;
  wire       [7:0]    _zz_invMixed_10_10;
  wire       [7:0]    _zz_invMixed_10_11;
  wire       [7:0]    _zz_invMixed_10_12;
  wire       [7:0]    _zz_invMixed_10_13;
  wire       [7:0]    _zz_invMixed_10_14;
  wire       [7:0]    _zz_invMixed_10_15;
  wire       [7:0]    _zz_invMixed_10_16;
  wire       [7:0]    _zz_invMixed_10_17;
  wire       [7:0]    _zz_invMixed_10_18;
  wire       [7:0]    _zz_invMixed_10_19;
  wire       [7:0]    _zz_invMixed_10_20;
  wire       [7:0]    _zz_invMixed_10_21;
  wire       [7:0]    _zz_invMixed_10_22;
  wire       [7:0]    _zz_invMixed_10_23;
  wire       [7:0]    _zz_invMixed_10_24;
  wire       [7:0]    _zz_invMixed_10_25;
  wire       [7:0]    _zz_invMixed_10_26;
  wire       [7:0]    _zz_invMixed_10_27;
  wire       [7:0]    _zz_invMixed_11;
  wire       [7:0]    _zz_invMixed_11_1;
  wire       [7:0]    _zz_invMixed_11_2;
  wire       [7:0]    _zz_invMixed_11_3;
  wire       [7:0]    _zz_invMixed_11_4;
  wire       [7:0]    _zz_invMixed_11_5;
  wire       [7:0]    _zz_invMixed_11_6;
  wire       [7:0]    _zz_invMixed_11_7;
  wire       [7:0]    _zz_invMixed_11_8;
  wire       [7:0]    _zz_invMixed_11_9;
  wire       [7:0]    _zz_invMixed_11_10;
  wire       [7:0]    _zz_invMixed_11_11;
  wire       [7:0]    _zz_invMixed_11_12;
  wire       [7:0]    _zz_invMixed_11_13;
  wire       [7:0]    _zz_invMixed_11_14;
  wire       [7:0]    _zz_invMixed_11_15;
  wire       [7:0]    _zz_invMixed_11_16;
  wire       [7:0]    _zz_invMixed_11_17;
  wire       [7:0]    _zz_invMixed_11_18;
  wire       [7:0]    _zz_invMixed_11_19;
  wire       [7:0]    _zz_invMixed_11_20;
  wire       [7:0]    _zz_invMixed_11_21;
  wire       [7:0]    _zz_invMixed_11_22;
  wire       [7:0]    _zz_invMixed_11_23;
  wire       [7:0]    _zz_invMixed_11_24;
  wire       [7:0]    _zz_invMixed_11_25;
  wire       [7:0]    _zz_invMixed_11_26;
  wire       [7:0]    _zz_invMixed_11_27;
  wire       [7:0]    _zz_invMixed_12_4;
  wire       [7:0]    _zz_invMixed_12_5;
  wire       [7:0]    _zz_invMixed_12_6;
  wire       [7:0]    _zz_invMixed_12_7;
  wire       [7:0]    _zz_invMixed_12_8;
  wire       [7:0]    _zz_invMixed_12_9;
  wire       [7:0]    _zz_invMixed_12_10;
  wire       [7:0]    _zz_invMixed_12_11;
  wire       [7:0]    _zz_invMixed_12_12;
  wire       [7:0]    _zz_invMixed_12_13;
  wire       [7:0]    _zz_invMixed_12_14;
  wire       [7:0]    _zz_invMixed_12_15;
  wire       [7:0]    _zz_invMixed_12_16;
  wire       [7:0]    _zz_invMixed_12_17;
  wire       [7:0]    _zz_invMixed_12_18;
  wire       [7:0]    _zz_invMixed_12_19;
  wire       [7:0]    _zz_invMixed_12_20;
  wire       [7:0]    _zz_invMixed_12_21;
  wire       [7:0]    _zz_invMixed_12_22;
  wire       [7:0]    _zz_invMixed_12_23;
  wire       [7:0]    _zz_invMixed_12_24;
  wire       [7:0]    _zz_invMixed_12_25;
  wire       [7:0]    _zz_invMixed_12_26;
  wire       [7:0]    _zz_invMixed_12_27;
  wire       [7:0]    _zz_invMixed_12_28;
  wire       [7:0]    _zz_invMixed_12_29;
  wire       [7:0]    _zz_invMixed_12_30;
  wire       [7:0]    _zz_invMixed_12_31;
  wire       [7:0]    _zz_invMixed_13;
  wire       [7:0]    _zz_invMixed_13_1;
  wire       [7:0]    _zz_invMixed_13_2;
  wire       [7:0]    _zz_invMixed_13_3;
  wire       [7:0]    _zz_invMixed_13_4;
  wire       [7:0]    _zz_invMixed_13_5;
  wire       [7:0]    _zz_invMixed_13_6;
  wire       [7:0]    _zz_invMixed_13_7;
  wire       [7:0]    _zz_invMixed_13_8;
  wire       [7:0]    _zz_invMixed_13_9;
  wire       [7:0]    _zz_invMixed_13_10;
  wire       [7:0]    _zz_invMixed_13_11;
  wire       [7:0]    _zz_invMixed_13_12;
  wire       [7:0]    _zz_invMixed_13_13;
  wire       [7:0]    _zz_invMixed_13_14;
  wire       [7:0]    _zz_invMixed_13_15;
  wire       [7:0]    _zz_invMixed_13_16;
  wire       [7:0]    _zz_invMixed_13_17;
  wire       [7:0]    _zz_invMixed_13_18;
  wire       [7:0]    _zz_invMixed_13_19;
  wire       [7:0]    _zz_invMixed_13_20;
  wire       [7:0]    _zz_invMixed_13_21;
  wire       [7:0]    _zz_invMixed_13_22;
  wire       [7:0]    _zz_invMixed_13_23;
  wire       [7:0]    _zz_invMixed_13_24;
  wire       [7:0]    _zz_invMixed_13_25;
  wire       [7:0]    _zz_invMixed_13_26;
  wire       [7:0]    _zz_invMixed_13_27;
  wire       [7:0]    _zz_invMixed_14;
  wire       [7:0]    _zz_invMixed_14_1;
  wire       [7:0]    _zz_invMixed_14_2;
  wire       [7:0]    _zz_invMixed_14_3;
  wire       [7:0]    _zz_invMixed_14_4;
  wire       [7:0]    _zz_invMixed_14_5;
  wire       [7:0]    _zz_invMixed_14_6;
  wire       [7:0]    _zz_invMixed_14_7;
  wire       [7:0]    _zz_invMixed_14_8;
  wire       [7:0]    _zz_invMixed_14_9;
  wire       [7:0]    _zz_invMixed_14_10;
  wire       [7:0]    _zz_invMixed_14_11;
  wire       [7:0]    _zz_invMixed_14_12;
  wire       [7:0]    _zz_invMixed_14_13;
  wire       [7:0]    _zz_invMixed_14_14;
  wire       [7:0]    _zz_invMixed_14_15;
  wire       [7:0]    _zz_invMixed_14_16;
  wire       [7:0]    _zz_invMixed_14_17;
  wire       [7:0]    _zz_invMixed_14_18;
  wire       [7:0]    _zz_invMixed_14_19;
  wire       [7:0]    _zz_invMixed_14_20;
  wire       [7:0]    _zz_invMixed_14_21;
  wire       [7:0]    _zz_invMixed_14_22;
  wire       [7:0]    _zz_invMixed_14_23;
  wire       [7:0]    _zz_invMixed_14_24;
  wire       [7:0]    _zz_invMixed_14_25;
  wire       [7:0]    _zz_invMixed_14_26;
  wire       [7:0]    _zz_invMixed_14_27;
  wire       [7:0]    _zz_invMixed_15;
  wire       [7:0]    _zz_invMixed_15_1;
  wire       [7:0]    _zz_invMixed_15_2;
  wire       [7:0]    _zz_invMixed_15_3;
  wire       [7:0]    _zz_invMixed_15_4;
  wire       [7:0]    _zz_invMixed_15_5;
  wire       [7:0]    _zz_invMixed_15_6;
  wire       [7:0]    _zz_invMixed_15_7;
  wire       [7:0]    _zz_invMixed_15_8;
  wire       [7:0]    _zz_invMixed_15_9;
  wire       [7:0]    _zz_invMixed_15_10;
  wire       [7:0]    _zz_invMixed_15_11;
  wire       [7:0]    _zz_invMixed_15_12;
  wire       [7:0]    _zz_invMixed_15_13;
  wire       [7:0]    _zz_invMixed_15_14;
  wire       [7:0]    _zz_invMixed_15_15;
  wire       [7:0]    _zz_invMixed_15_16;
  wire       [7:0]    _zz_invMixed_15_17;
  wire       [7:0]    _zz_invMixed_15_18;
  wire       [7:0]    _zz_invMixed_15_19;
  wire       [7:0]    _zz_invMixed_15_20;
  wire       [7:0]    _zz_invMixed_15_21;
  wire       [7:0]    _zz_invMixed_15_22;
  wire       [7:0]    _zz_invMixed_15_23;
  wire       [7:0]    _zz_invMixed_15_24;
  wire       [7:0]    _zz_invMixed_15_25;
  wire       [7:0]    _zz_invMixed_15_26;
  wire       [7:0]    _zz_invMixed_15_27;
  wire                when_AES128_l397;
  wire                when_AES128_l403;
  wire                when_AES128_l244;
  wire                when_AES128_l315;
  wire                when_AES128_l339;

  assign _zz__zz_stateReg_36 = ({1'd0,_zz_stateReg_4} <<< 1'd1);
  assign _zz__zz_stateReg_37 = ({1'd0,_zz_stateReg_5} <<< 1'd1);
  assign _zz__zz_stateReg_38 = ({1'd0,_zz_stateReg_5} <<< 1'd1);
  assign _zz__zz_stateReg_39 = ({1'd0,_zz_stateReg_6} <<< 1'd1);
  assign _zz__zz_stateReg_40 = ({1'd0,_zz_stateReg_6} <<< 1'd1);
  assign _zz__zz_stateReg_41 = ({1'd0,_zz_stateReg_7} <<< 1'd1);
  assign _zz__zz_stateReg_42 = ({1'd0,_zz_stateReg_4} <<< 1'd1);
  assign _zz__zz_stateReg_43 = ({1'd0,_zz_stateReg_7} <<< 1'd1);
  assign _zz__zz_stateReg_44 = ({1'd0,_zz_stateReg_8} <<< 1'd1);
  assign _zz__zz_stateReg_45 = ({1'd0,_zz_stateReg_9} <<< 1'd1);
  assign _zz__zz_stateReg_46 = ({1'd0,_zz_stateReg_9} <<< 1'd1);
  assign _zz__zz_stateReg_47 = ({1'd0,_zz_stateReg_10} <<< 1'd1);
  assign _zz__zz_stateReg_48 = ({1'd0,_zz_stateReg_10} <<< 1'd1);
  assign _zz__zz_stateReg_49 = ({1'd0,_zz_stateReg_11} <<< 1'd1);
  assign _zz__zz_stateReg_50 = ({1'd0,_zz_stateReg_8} <<< 1'd1);
  assign _zz__zz_stateReg_51 = ({1'd0,_zz_stateReg_11} <<< 1'd1);
  assign _zz__zz_stateReg_52 = ({1'd0,_zz_stateReg_12} <<< 1'd1);
  assign _zz__zz_stateReg_53 = ({1'd0,_zz_stateReg_13} <<< 1'd1);
  assign _zz__zz_stateReg_54 = ({1'd0,_zz_stateReg_13} <<< 1'd1);
  assign _zz__zz_stateReg_55 = ({1'd0,_zz_stateReg_14} <<< 1'd1);
  assign _zz__zz_stateReg_56 = ({1'd0,_zz_stateReg_14} <<< 1'd1);
  assign _zz__zz_stateReg_57 = ({1'd0,_zz_stateReg_15} <<< 1'd1);
  assign _zz__zz_stateReg_58 = ({1'd0,_zz_stateReg_12} <<< 1'd1);
  assign _zz__zz_stateReg_59 = ({1'd0,_zz_stateReg_15} <<< 1'd1);
  assign _zz__zz_stateReg_60 = ({1'd0,_zz_stateReg_16} <<< 1'd1);
  assign _zz__zz_stateReg_61 = ({1'd0,_zz_stateReg_17} <<< 1'd1);
  assign _zz__zz_stateReg_62 = ({1'd0,_zz_stateReg_17} <<< 1'd1);
  assign _zz__zz_stateReg_63 = ({1'd0,_zz_stateReg_18} <<< 1'd1);
  assign _zz__zz_stateReg_64 = ({1'd0,_zz_stateReg_18} <<< 1'd1);
  assign _zz__zz_stateReg_65 = ({1'd0,_zz_stateReg_19} <<< 1'd1);
  assign _zz__zz_stateReg_66 = ({1'd0,_zz_stateReg_16} <<< 1'd1);
  assign _zz__zz_stateReg_67 = ({1'd0,_zz_stateReg_19} <<< 1'd1);
  assign _zz__zz_invMixed_0_5_1 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_0_7_1 = ({1'd0,_zz_invMixed_0_6} <<< 1'd1);
  assign _zz__zz_invMixed_0_9_1 = ({1'd0,_zz_invMixed_0_8} <<< 1'd1);
  assign _zz__zz_invMixed_0_10_1 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_0_12_1 = ({1'd0,_zz_invMixed_0_11} <<< 1'd1);
  assign _zz__zz_invMixed_0_13_1 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_0_14_1 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_0_16 = ({1'd0,_zz_invMixed_0_15} <<< 1'd1);
  assign _zz__zz_invMixed_0_18 = ({1'd0,_zz_invMixed_0_17} <<< 1'd1);
  assign _zz__zz_invMixed_0_19 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_0_20 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_0_22 = ({1'd0,_zz_invMixed_0_21} <<< 1'd1);
  assign _zz__zz_invMixed_0_24 = ({1'd0,_zz_invMixed_0_23} <<< 1'd1);
  assign _zz__zz_invMixed_0_25 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_0_27 = ({1'd0,_zz_invMixed_0_26} <<< 1'd1);
  assign _zz__zz_invMixed_0_28 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_0_30 = ({1'd0,_zz_invMixed_0_29} <<< 1'd1);
  assign _zz__zz_invMixed_0_32 = ({1'd0,_zz_invMixed_0_31} <<< 1'd1);
  assign _zz__zz_invMixed_1 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_1_2 = ({1'd0,_zz_invMixed_1_1} <<< 1'd1);
  assign _zz__zz_invMixed_1_4 = ({1'd0,_zz_invMixed_1_3} <<< 1'd1);
  assign _zz__zz_invMixed_1_5 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_1_7 = ({1'd0,_zz_invMixed_1_6} <<< 1'd1);
  assign _zz__zz_invMixed_1_9 = ({1'd0,_zz_invMixed_1_8} <<< 1'd1);
  assign _zz__zz_invMixed_1_10 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_1_12 = ({1'd0,_zz_invMixed_1_11} <<< 1'd1);
  assign _zz__zz_invMixed_1_13 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_1_14 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_1_16 = ({1'd0,_zz_invMixed_1_15} <<< 1'd1);
  assign _zz__zz_invMixed_1_18 = ({1'd0,_zz_invMixed_1_17} <<< 1'd1);
  assign _zz__zz_invMixed_1_19 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_1_20 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_1_22 = ({1'd0,_zz_invMixed_1_21} <<< 1'd1);
  assign _zz__zz_invMixed_1_24 = ({1'd0,_zz_invMixed_1_23} <<< 1'd1);
  assign _zz__zz_invMixed_1_25 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_1_27 = ({1'd0,_zz_invMixed_1_26} <<< 1'd1);
  assign _zz__zz_invMixed_2 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_2_2 = ({1'd0,_zz_invMixed_2_1} <<< 1'd1);
  assign _zz__zz_invMixed_2_4 = ({1'd0,_zz_invMixed_2_3} <<< 1'd1);
  assign _zz__zz_invMixed_2_5 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_2_7 = ({1'd0,_zz_invMixed_2_6} <<< 1'd1);
  assign _zz__zz_invMixed_2_8 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_2_10 = ({1'd0,_zz_invMixed_2_9} <<< 1'd1);
  assign _zz__zz_invMixed_2_12 = ({1'd0,_zz_invMixed_2_11} <<< 1'd1);
  assign _zz__zz_invMixed_2_13 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_2_15 = ({1'd0,_zz_invMixed_2_14} <<< 1'd1);
  assign _zz__zz_invMixed_2_17 = ({1'd0,_zz_invMixed_2_16} <<< 1'd1);
  assign _zz__zz_invMixed_2_18 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_2_20 = ({1'd0,_zz_invMixed_2_19} <<< 1'd1);
  assign _zz__zz_invMixed_2_21 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_2_22 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_2_24 = ({1'd0,_zz_invMixed_2_23} <<< 1'd1);
  assign _zz__zz_invMixed_2_26 = ({1'd0,_zz_invMixed_2_25} <<< 1'd1);
  assign _zz__zz_invMixed_2_27 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_3 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_3_2 = ({1'd0,_zz_invMixed_3_1} <<< 1'd1);
  assign _zz__zz_invMixed_3_4 = ({1'd0,_zz_invMixed_3_3} <<< 1'd1);
  assign _zz__zz_invMixed_3_5 = ({1'd0,_zz_invMixed_0_1} <<< 1'd1);
  assign _zz__zz_invMixed_3_6 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_3_8 = ({1'd0,_zz_invMixed_3_7} <<< 1'd1);
  assign _zz__zz_invMixed_3_10 = ({1'd0,_zz_invMixed_3_9} <<< 1'd1);
  assign _zz__zz_invMixed_3_11 = ({1'd0,_zz_invMixed_0_2} <<< 1'd1);
  assign _zz__zz_invMixed_3_13 = ({1'd0,_zz_invMixed_3_12} <<< 1'd1);
  assign _zz__zz_invMixed_3_14 = ({1'd0,_zz_invMixed_0_3} <<< 1'd1);
  assign _zz__zz_invMixed_3_16 = ({1'd0,_zz_invMixed_3_15} <<< 1'd1);
  assign _zz__zz_invMixed_3_18 = ({1'd0,_zz_invMixed_3_17} <<< 1'd1);
  assign _zz__zz_invMixed_3_19 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_3_21 = ({1'd0,_zz_invMixed_3_20} <<< 1'd1);
  assign _zz__zz_invMixed_3_23 = ({1'd0,_zz_invMixed_3_22} <<< 1'd1);
  assign _zz__zz_invMixed_3_24 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_3_26 = ({1'd0,_zz_invMixed_3_25} <<< 1'd1);
  assign _zz__zz_invMixed_3_27 = ({1'd0,_zz_invMixed_0_4} <<< 1'd1);
  assign _zz__zz_invMixed_4_4 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_4_6 = ({1'd0,_zz_invMixed_4_5} <<< 1'd1);
  assign _zz__zz_invMixed_4_8 = ({1'd0,_zz_invMixed_4_7} <<< 1'd1);
  assign _zz__zz_invMixed_4_9 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_4_11 = ({1'd0,_zz_invMixed_4_10} <<< 1'd1);
  assign _zz__zz_invMixed_4_12 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_4_13 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_4_15 = ({1'd0,_zz_invMixed_4_14} <<< 1'd1);
  assign _zz__zz_invMixed_4_17 = ({1'd0,_zz_invMixed_4_16} <<< 1'd1);
  assign _zz__zz_invMixed_4_18 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_4_19 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_4_21 = ({1'd0,_zz_invMixed_4_20} <<< 1'd1);
  assign _zz__zz_invMixed_4_23 = ({1'd0,_zz_invMixed_4_22} <<< 1'd1);
  assign _zz__zz_invMixed_4_24 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_4_26 = ({1'd0,_zz_invMixed_4_25} <<< 1'd1);
  assign _zz__zz_invMixed_4_27 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_4_29 = ({1'd0,_zz_invMixed_4_28} <<< 1'd1);
  assign _zz__zz_invMixed_4_31 = ({1'd0,_zz_invMixed_4_30} <<< 1'd1);
  assign _zz__zz_invMixed_5 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_5_2 = ({1'd0,_zz_invMixed_5_1} <<< 1'd1);
  assign _zz__zz_invMixed_5_4 = ({1'd0,_zz_invMixed_5_3} <<< 1'd1);
  assign _zz__zz_invMixed_5_5 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_5_7 = ({1'd0,_zz_invMixed_5_6} <<< 1'd1);
  assign _zz__zz_invMixed_5_9 = ({1'd0,_zz_invMixed_5_8} <<< 1'd1);
  assign _zz__zz_invMixed_5_10 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_5_12 = ({1'd0,_zz_invMixed_5_11} <<< 1'd1);
  assign _zz__zz_invMixed_5_13 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_5_14 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_5_16 = ({1'd0,_zz_invMixed_5_15} <<< 1'd1);
  assign _zz__zz_invMixed_5_18 = ({1'd0,_zz_invMixed_5_17} <<< 1'd1);
  assign _zz__zz_invMixed_5_19 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_5_20 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_5_22 = ({1'd0,_zz_invMixed_5_21} <<< 1'd1);
  assign _zz__zz_invMixed_5_24 = ({1'd0,_zz_invMixed_5_23} <<< 1'd1);
  assign _zz__zz_invMixed_5_25 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_5_27 = ({1'd0,_zz_invMixed_5_26} <<< 1'd1);
  assign _zz__zz_invMixed_6 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_6_2 = ({1'd0,_zz_invMixed_6_1} <<< 1'd1);
  assign _zz__zz_invMixed_6_4 = ({1'd0,_zz_invMixed_6_3} <<< 1'd1);
  assign _zz__zz_invMixed_6_5 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_6_7 = ({1'd0,_zz_invMixed_6_6} <<< 1'd1);
  assign _zz__zz_invMixed_6_8 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_6_10 = ({1'd0,_zz_invMixed_6_9} <<< 1'd1);
  assign _zz__zz_invMixed_6_12 = ({1'd0,_zz_invMixed_6_11} <<< 1'd1);
  assign _zz__zz_invMixed_6_13 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_6_15 = ({1'd0,_zz_invMixed_6_14} <<< 1'd1);
  assign _zz__zz_invMixed_6_17 = ({1'd0,_zz_invMixed_6_16} <<< 1'd1);
  assign _zz__zz_invMixed_6_18 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_6_20 = ({1'd0,_zz_invMixed_6_19} <<< 1'd1);
  assign _zz__zz_invMixed_6_21 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_6_22 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_6_24 = ({1'd0,_zz_invMixed_6_23} <<< 1'd1);
  assign _zz__zz_invMixed_6_26 = ({1'd0,_zz_invMixed_6_25} <<< 1'd1);
  assign _zz__zz_invMixed_6_27 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_7 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_7_2 = ({1'd0,_zz_invMixed_7_1} <<< 1'd1);
  assign _zz__zz_invMixed_7_4 = ({1'd0,_zz_invMixed_7_3} <<< 1'd1);
  assign _zz__zz_invMixed_7_5 = ({1'd0,_zz_invMixed_4} <<< 1'd1);
  assign _zz__zz_invMixed_7_6 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_7_8 = ({1'd0,_zz_invMixed_7_7} <<< 1'd1);
  assign _zz__zz_invMixed_7_10 = ({1'd0,_zz_invMixed_7_9} <<< 1'd1);
  assign _zz__zz_invMixed_7_11 = ({1'd0,_zz_invMixed_4_1} <<< 1'd1);
  assign _zz__zz_invMixed_7_13 = ({1'd0,_zz_invMixed_7_12} <<< 1'd1);
  assign _zz__zz_invMixed_7_14 = ({1'd0,_zz_invMixed_4_2} <<< 1'd1);
  assign _zz__zz_invMixed_7_16 = ({1'd0,_zz_invMixed_7_15} <<< 1'd1);
  assign _zz__zz_invMixed_7_18 = ({1'd0,_zz_invMixed_7_17} <<< 1'd1);
  assign _zz__zz_invMixed_7_19 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_7_21 = ({1'd0,_zz_invMixed_7_20} <<< 1'd1);
  assign _zz__zz_invMixed_7_23 = ({1'd0,_zz_invMixed_7_22} <<< 1'd1);
  assign _zz__zz_invMixed_7_24 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_7_26 = ({1'd0,_zz_invMixed_7_25} <<< 1'd1);
  assign _zz__zz_invMixed_7_27 = ({1'd0,_zz_invMixed_4_3} <<< 1'd1);
  assign _zz__zz_invMixed_8_4 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_8_6 = ({1'd0,_zz_invMixed_8_5} <<< 1'd1);
  assign _zz__zz_invMixed_8_8 = ({1'd0,_zz_invMixed_8_7} <<< 1'd1);
  assign _zz__zz_invMixed_8_9 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_8_11 = ({1'd0,_zz_invMixed_8_10} <<< 1'd1);
  assign _zz__zz_invMixed_8_12 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_8_13 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_8_15 = ({1'd0,_zz_invMixed_8_14} <<< 1'd1);
  assign _zz__zz_invMixed_8_17 = ({1'd0,_zz_invMixed_8_16} <<< 1'd1);
  assign _zz__zz_invMixed_8_18 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_8_19 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_8_21 = ({1'd0,_zz_invMixed_8_20} <<< 1'd1);
  assign _zz__zz_invMixed_8_23 = ({1'd0,_zz_invMixed_8_22} <<< 1'd1);
  assign _zz__zz_invMixed_8_24 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_8_26 = ({1'd0,_zz_invMixed_8_25} <<< 1'd1);
  assign _zz__zz_invMixed_8_27 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_8_29 = ({1'd0,_zz_invMixed_8_28} <<< 1'd1);
  assign _zz__zz_invMixed_8_31 = ({1'd0,_zz_invMixed_8_30} <<< 1'd1);
  assign _zz__zz_invMixed_9 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_9_2 = ({1'd0,_zz_invMixed_9_1} <<< 1'd1);
  assign _zz__zz_invMixed_9_4 = ({1'd0,_zz_invMixed_9_3} <<< 1'd1);
  assign _zz__zz_invMixed_9_5 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_9_7 = ({1'd0,_zz_invMixed_9_6} <<< 1'd1);
  assign _zz__zz_invMixed_9_9 = ({1'd0,_zz_invMixed_9_8} <<< 1'd1);
  assign _zz__zz_invMixed_9_10 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_9_12 = ({1'd0,_zz_invMixed_9_11} <<< 1'd1);
  assign _zz__zz_invMixed_9_13 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_9_14 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_9_16 = ({1'd0,_zz_invMixed_9_15} <<< 1'd1);
  assign _zz__zz_invMixed_9_18 = ({1'd0,_zz_invMixed_9_17} <<< 1'd1);
  assign _zz__zz_invMixed_9_19 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_9_20 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_9_22 = ({1'd0,_zz_invMixed_9_21} <<< 1'd1);
  assign _zz__zz_invMixed_9_24 = ({1'd0,_zz_invMixed_9_23} <<< 1'd1);
  assign _zz__zz_invMixed_9_25 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_9_27 = ({1'd0,_zz_invMixed_9_26} <<< 1'd1);
  assign _zz__zz_invMixed_10 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_10_2 = ({1'd0,_zz_invMixed_10_1} <<< 1'd1);
  assign _zz__zz_invMixed_10_4 = ({1'd0,_zz_invMixed_10_3} <<< 1'd1);
  assign _zz__zz_invMixed_10_5 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_10_7 = ({1'd0,_zz_invMixed_10_6} <<< 1'd1);
  assign _zz__zz_invMixed_10_8 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_10_10 = ({1'd0,_zz_invMixed_10_9} <<< 1'd1);
  assign _zz__zz_invMixed_10_12 = ({1'd0,_zz_invMixed_10_11} <<< 1'd1);
  assign _zz__zz_invMixed_10_13 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_10_15 = ({1'd0,_zz_invMixed_10_14} <<< 1'd1);
  assign _zz__zz_invMixed_10_17 = ({1'd0,_zz_invMixed_10_16} <<< 1'd1);
  assign _zz__zz_invMixed_10_18 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_10_20 = ({1'd0,_zz_invMixed_10_19} <<< 1'd1);
  assign _zz__zz_invMixed_10_21 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_10_22 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_10_24 = ({1'd0,_zz_invMixed_10_23} <<< 1'd1);
  assign _zz__zz_invMixed_10_26 = ({1'd0,_zz_invMixed_10_25} <<< 1'd1);
  assign _zz__zz_invMixed_10_27 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_11 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_11_2 = ({1'd0,_zz_invMixed_11_1} <<< 1'd1);
  assign _zz__zz_invMixed_11_4 = ({1'd0,_zz_invMixed_11_3} <<< 1'd1);
  assign _zz__zz_invMixed_11_5 = ({1'd0,_zz_invMixed_8} <<< 1'd1);
  assign _zz__zz_invMixed_11_6 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_11_8 = ({1'd0,_zz_invMixed_11_7} <<< 1'd1);
  assign _zz__zz_invMixed_11_10 = ({1'd0,_zz_invMixed_11_9} <<< 1'd1);
  assign _zz__zz_invMixed_11_11 = ({1'd0,_zz_invMixed_8_1} <<< 1'd1);
  assign _zz__zz_invMixed_11_13 = ({1'd0,_zz_invMixed_11_12} <<< 1'd1);
  assign _zz__zz_invMixed_11_14 = ({1'd0,_zz_invMixed_8_2} <<< 1'd1);
  assign _zz__zz_invMixed_11_16 = ({1'd0,_zz_invMixed_11_15} <<< 1'd1);
  assign _zz__zz_invMixed_11_18 = ({1'd0,_zz_invMixed_11_17} <<< 1'd1);
  assign _zz__zz_invMixed_11_19 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_11_21 = ({1'd0,_zz_invMixed_11_20} <<< 1'd1);
  assign _zz__zz_invMixed_11_23 = ({1'd0,_zz_invMixed_11_22} <<< 1'd1);
  assign _zz__zz_invMixed_11_24 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_11_26 = ({1'd0,_zz_invMixed_11_25} <<< 1'd1);
  assign _zz__zz_invMixed_11_27 = ({1'd0,_zz_invMixed_8_3} <<< 1'd1);
  assign _zz__zz_invMixed_12_4 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_12_6 = ({1'd0,_zz_invMixed_12_5} <<< 1'd1);
  assign _zz__zz_invMixed_12_8 = ({1'd0,_zz_invMixed_12_7} <<< 1'd1);
  assign _zz__zz_invMixed_12_9 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_12_11 = ({1'd0,_zz_invMixed_12_10} <<< 1'd1);
  assign _zz__zz_invMixed_12_12 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_12_13 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_12_15 = ({1'd0,_zz_invMixed_12_14} <<< 1'd1);
  assign _zz__zz_invMixed_12_17 = ({1'd0,_zz_invMixed_12_16} <<< 1'd1);
  assign _zz__zz_invMixed_12_18 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_12_19 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_12_21 = ({1'd0,_zz_invMixed_12_20} <<< 1'd1);
  assign _zz__zz_invMixed_12_23 = ({1'd0,_zz_invMixed_12_22} <<< 1'd1);
  assign _zz__zz_invMixed_12_24 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_12_26 = ({1'd0,_zz_invMixed_12_25} <<< 1'd1);
  assign _zz__zz_invMixed_12_27 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_12_29 = ({1'd0,_zz_invMixed_12_28} <<< 1'd1);
  assign _zz__zz_invMixed_12_31 = ({1'd0,_zz_invMixed_12_30} <<< 1'd1);
  assign _zz__zz_invMixed_13 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_13_2 = ({1'd0,_zz_invMixed_13_1} <<< 1'd1);
  assign _zz__zz_invMixed_13_4 = ({1'd0,_zz_invMixed_13_3} <<< 1'd1);
  assign _zz__zz_invMixed_13_5 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_13_7 = ({1'd0,_zz_invMixed_13_6} <<< 1'd1);
  assign _zz__zz_invMixed_13_9 = ({1'd0,_zz_invMixed_13_8} <<< 1'd1);
  assign _zz__zz_invMixed_13_10 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_13_12 = ({1'd0,_zz_invMixed_13_11} <<< 1'd1);
  assign _zz__zz_invMixed_13_13 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_13_14 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_13_16 = ({1'd0,_zz_invMixed_13_15} <<< 1'd1);
  assign _zz__zz_invMixed_13_18 = ({1'd0,_zz_invMixed_13_17} <<< 1'd1);
  assign _zz__zz_invMixed_13_19 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_13_20 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_13_22 = ({1'd0,_zz_invMixed_13_21} <<< 1'd1);
  assign _zz__zz_invMixed_13_24 = ({1'd0,_zz_invMixed_13_23} <<< 1'd1);
  assign _zz__zz_invMixed_13_25 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_13_27 = ({1'd0,_zz_invMixed_13_26} <<< 1'd1);
  assign _zz__zz_invMixed_14 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_14_2 = ({1'd0,_zz_invMixed_14_1} <<< 1'd1);
  assign _zz__zz_invMixed_14_4 = ({1'd0,_zz_invMixed_14_3} <<< 1'd1);
  assign _zz__zz_invMixed_14_5 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_14_7 = ({1'd0,_zz_invMixed_14_6} <<< 1'd1);
  assign _zz__zz_invMixed_14_8 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_14_10 = ({1'd0,_zz_invMixed_14_9} <<< 1'd1);
  assign _zz__zz_invMixed_14_12 = ({1'd0,_zz_invMixed_14_11} <<< 1'd1);
  assign _zz__zz_invMixed_14_13 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_14_15 = ({1'd0,_zz_invMixed_14_14} <<< 1'd1);
  assign _zz__zz_invMixed_14_17 = ({1'd0,_zz_invMixed_14_16} <<< 1'd1);
  assign _zz__zz_invMixed_14_18 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_14_20 = ({1'd0,_zz_invMixed_14_19} <<< 1'd1);
  assign _zz__zz_invMixed_14_21 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_14_22 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_14_24 = ({1'd0,_zz_invMixed_14_23} <<< 1'd1);
  assign _zz__zz_invMixed_14_26 = ({1'd0,_zz_invMixed_14_25} <<< 1'd1);
  assign _zz__zz_invMixed_14_27 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_15 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_15_2 = ({1'd0,_zz_invMixed_15_1} <<< 1'd1);
  assign _zz__zz_invMixed_15_4 = ({1'd0,_zz_invMixed_15_3} <<< 1'd1);
  assign _zz__zz_invMixed_15_5 = ({1'd0,_zz_invMixed_12} <<< 1'd1);
  assign _zz__zz_invMixed_15_6 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_15_8 = ({1'd0,_zz_invMixed_15_7} <<< 1'd1);
  assign _zz__zz_invMixed_15_10 = ({1'd0,_zz_invMixed_15_9} <<< 1'd1);
  assign _zz__zz_invMixed_15_11 = ({1'd0,_zz_invMixed_12_1} <<< 1'd1);
  assign _zz__zz_invMixed_15_13 = ({1'd0,_zz_invMixed_15_12} <<< 1'd1);
  assign _zz__zz_invMixed_15_14 = ({1'd0,_zz_invMixed_12_2} <<< 1'd1);
  assign _zz__zz_invMixed_15_16 = ({1'd0,_zz_invMixed_15_15} <<< 1'd1);
  assign _zz__zz_invMixed_15_18 = ({1'd0,_zz_invMixed_15_17} <<< 1'd1);
  assign _zz__zz_invMixed_15_19 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_15_21 = ({1'd0,_zz_invMixed_15_20} <<< 1'd1);
  assign _zz__zz_invMixed_15_23 = ({1'd0,_zz_invMixed_15_22} <<< 1'd1);
  assign _zz__zz_invMixed_15_24 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_invMixed_15_26 = ({1'd0,_zz_invMixed_15_25} <<< 1'd1);
  assign _zz__zz_invMixed_15_27 = ({1'd0,_zz_invMixed_12_3} <<< 1'd1);
  assign _zz__zz_stateReg_4_1 = stateReg[127 : 120];
  assign _zz__zz_stateReg_8_1 = stateReg[95 : 88];
  assign _zz__zz_stateReg_12_1 = stateReg[63 : 56];
  assign _zz__zz_stateReg_16_1 = stateReg[31 : 24];
  assign _zz__zz_stateReg_5_1 = stateReg[87 : 80];
  assign _zz__zz_stateReg_9_1 = stateReg[55 : 48];
  assign _zz__zz_stateReg_13_1 = stateReg[23 : 16];
  assign _zz__zz_stateReg_17_1 = stateReg[119 : 112];
  assign _zz__zz_stateReg_6_1 = stateReg[47 : 40];
  assign _zz__zz_stateReg_10_1 = stateReg[15 : 8];
  assign _zz__zz_stateReg_14_1 = stateReg[111 : 104];
  assign _zz__zz_stateReg_18_1 = stateReg[79 : 72];
  assign _zz__zz_stateReg_7_1 = stateReg[7 : 0];
  assign _zz__zz_stateReg_11_1 = stateReg[103 : 96];
  assign _zz__zz_stateReg_15_1 = stateReg[71 : 64];
  assign _zz__zz_stateReg_19_1 = stateReg[39 : 32];
  assign _zz__zz_roundKeyReg_0_2_1 = _zz_roundKeyReg_0_1[31 : 24];
  assign _zz__zz_roundKeyReg_0_2_3 = _zz_roundKeyReg_0_1[23 : 16];
  assign _zz__zz_roundKeyReg_0_2_5 = _zz_roundKeyReg_0_1[15 : 8];
  assign _zz__zz_roundKeyReg_0_2_7 = _zz_roundKeyReg_0_1[7 : 0];
  assign _zz__zz_stateReg_71_1 = _zz_stateReg_70[31 : 24];
  assign _zz__zz_stateReg_71_3 = _zz_stateReg_70[23 : 16];
  assign _zz__zz_stateReg_71_5 = _zz_stateReg_70[15 : 8];
  assign _zz__zz_stateReg_71_7 = _zz_stateReg_70[7 : 0];
  assign _zz__zz_roundKeyReg_0_5_1 = _zz_roundKeyReg_0_4[31 : 24];
  assign _zz__zz_roundKeyReg_0_5_3 = _zz_roundKeyReg_0_4[23 : 16];
  assign _zz__zz_roundKeyReg_0_5_5 = _zz_roundKeyReg_0_4[15 : 8];
  assign _zz__zz_roundKeyReg_0_5_7 = _zz_roundKeyReg_0_4[7 : 0];
  assign _zz_stateReg_75 = {{{{{_zz_stateReg_76,_zz_stateReg_82},_zz_stateReg_83},(_zz_stateReg_84 ^ _zz_stateReg_85)},(_zz_stateReg_86 ^ _zz_stateReg_2[31 : 24])},(io_dataIn[55 : 48] ^ _zz_stateReg_2[23 : 16])};
  assign _zz_stateReg_87 = (io_dataIn[47 : 40] ^ _zz_stateReg_2[15 : 8]);
  assign _zz_stateReg_88 = (io_dataIn[39 : 32] ^ _zz_stateReg_2[7 : 0]);
  assign _zz_stateReg_89 = io_dataIn[31 : 24];
  assign _zz_stateReg_90 = _zz_stateReg_3[31 : 24];
  assign _zz_stateReg_91 = io_dataIn[23 : 16];
  assign _zz_stateReg_76 = {{{{_zz_stateReg_77,_zz_stateReg_78},(_zz_stateReg_79 ^ _zz_stateReg_80)},(_zz_stateReg_81 ^ _zz_stateReg[7 : 0])},(io_dataIn[95 : 88] ^ _zz_stateReg_1[31 : 24])};
  assign _zz_stateReg_82 = (io_dataIn[87 : 80] ^ _zz_stateReg_1[23 : 16]);
  assign _zz_stateReg_83 = (io_dataIn[79 : 72] ^ _zz_stateReg_1[15 : 8]);
  assign _zz_stateReg_84 = io_dataIn[71 : 64];
  assign _zz_stateReg_85 = _zz_stateReg_1[7 : 0];
  assign _zz_stateReg_86 = io_dataIn[63 : 56];
  assign _zz_stateReg_77 = (io_dataIn[127 : 120] ^ _zz_stateReg[31 : 24]);
  assign _zz_stateReg_78 = (io_dataIn[119 : 112] ^ _zz_stateReg[23 : 16]);
  assign _zz_stateReg_79 = io_dataIn[111 : 104];
  assign _zz_stateReg_80 = _zz_stateReg[15 : 8];
  assign _zz_stateReg_81 = io_dataIn[103 : 96];
  assign _zz__zz_stateReg_68 = {{{{_zz_stateReg_20,_zz_stateReg_21},_zz_stateReg_22},_zz_stateReg_23},_zz_stateReg_24};
  assign _zz__zz_stateReg_68_1 = _zz_stateReg_25;
  assign _zz__zz_stateReg_69 = {{{{{{_zz_roundKeyReg_0_2[31 : 24],_zz_roundKeyReg_0_2[23 : 16]},_zz_roundKeyReg_0_2[15 : 8]},_zz_roundKeyReg_0_2[7 : 0]},_zz_roundKeyReg_1[31 : 24]},_zz_roundKeyReg_1[23 : 16]},_zz_roundKeyReg_1[15 : 8]};
  assign _zz__zz_stateReg_69_1 = _zz_roundKeyReg_1[7 : 0];
  assign _zz__zz_stateReg_69_2 = _zz_roundKeyReg_2[31 : 24];
  assign _zz_stateReg_92 = {{{{{{_zz_stateReg_71[31 : 24],_zz_stateReg_71[23 : 16]},_zz_stateReg_71[15 : 8]},_zz_stateReg_71[7 : 0]},_zz_stateReg_72[31 : 24]},_zz_stateReg_72[23 : 16]},_zz_stateReg_72[15 : 8]};
  assign _zz_stateReg_93 = _zz_stateReg_72[7 : 0];
  assign _zz_stateReg_94 = _zz_stateReg_73[31 : 24];
  assign _zz__zz_invMixed_0 = {{{{{_zz__zz_invMixed_0_1,_zz__zz_invMixed_0_4},invSub_7},invSub_8},invSub_9},invSub_10};
  assign _zz__zz_invMixed_0_5 = invSub_11;
  assign _zz__zz_invMixed_0_6 = {{{{{_zz__zz_invMixed_0_7,_zz__zz_invMixed_0_11},_zz__zz_invMixed_0_12},_zz_roundKeyReg_2_2[31 : 24]},_zz_roundKeyReg_2_2[23 : 16]},_zz_roundKeyReg_2_2[15 : 8]};
  assign _zz__zz_invMixed_0_13 = _zz_roundKeyReg_2_2[7 : 0];
  assign _zz__zz_invMixed_0_14 = _zz_roundKeyReg_3_2[31 : 24];
  assign _zz__zz_invMixed_0_1 = {{{{{_zz__zz_invMixed_0_2,_zz__zz_invMixed_0_3},invSub_2},invSub_3},invSub_4},invSub_5};
  assign _zz__zz_invMixed_0_4 = invSub_6;
  assign _zz__zz_invMixed_0_7 = {{{{{_zz__zz_invMixed_0_8,_zz__zz_invMixed_0_9},_zz__zz_invMixed_0_10},_zz_roundKeyReg_0_5[7 : 0]},_zz_roundKeyReg_1_2[31 : 24]},_zz_roundKeyReg_1_2[23 : 16]};
  assign _zz__zz_invMixed_0_11 = _zz_roundKeyReg_1_2[15 : 8];
  assign _zz__zz_invMixed_0_12 = _zz_roundKeyReg_1_2[7 : 0];
  assign _zz__zz_invMixed_0_2 = invSub_0;
  assign _zz__zz_invMixed_0_3 = invSub_1;
  assign _zz__zz_invMixed_0_8 = _zz_roundKeyReg_0_5[31 : 24];
  assign _zz__zz_invMixed_0_9 = _zz_roundKeyReg_0_5[23 : 16];
  assign _zz__zz_invMixed_0_10 = _zz_roundKeyReg_0_5[15 : 8];
  assign _zz_invMixed_0_33 = (_zz_invMixed_0_8[7] ? (_zz_invMixed_0_9 ^ 8'h1b) : _zz_invMixed_0_9);
  assign _zz_invMixed_0_34 = (_zz_invMixed_0_11[7] ? (_zz_invMixed_0_12 ^ 8'h1b) : _zz_invMixed_0_12);
  assign _zz_invMixed_0_35 = _zz_invMixed_0_1[7];
  assign _zz_invMixed_0_36 = (_zz_invMixed_0_13 ^ 8'h1b);
  assign _zz_invMixed_0_37 = (_zz_invMixed_0_17[7] ? (_zz_invMixed_0_18 ^ 8'h1b) : _zz_invMixed_0_18);
  assign _zz_invMixed_0_38 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_0_19 ^ 8'h1b) : _zz_invMixed_0_19);
  assign _zz_invMixed_0_39 = _zz_invMixed_0_23[7];
  assign _zz_invMixed_0_40 = (_zz_invMixed_0_24 ^ 8'h1b);
  assign _zz_invMixed_0_41 = _zz_invMixed_0_26[7];
  assign _zz_invMixed_0_42 = (_zz_invMixed_0_27 ^ 8'h1b);
  assign _zz_invMixed_1_28 = _zz_invMixed_1_3[7];
  assign _zz_invMixed_1_29 = (_zz_invMixed_1_4 ^ 8'h1b);
  assign _zz_invMixed_1_30 = (_zz_invMixed_1_8[7] ? (_zz_invMixed_1_9 ^ 8'h1b) : _zz_invMixed_1_9);
  assign _zz_invMixed_1_31 = (_zz_invMixed_1_11[7] ? (_zz_invMixed_1_12 ^ 8'h1b) : _zz_invMixed_1_12);
  assign _zz_invMixed_1_32 = _zz_invMixed_0_2[7];
  assign _zz_invMixed_1_33 = (_zz_invMixed_1_13 ^ 8'h1b);
  assign _zz_invMixed_1_34 = _zz_invMixed_1_17[7];
  assign _zz_invMixed_1_35 = (_zz_invMixed_1_18 ^ 8'h1b);
  assign _zz_invMixed_1_36 = _zz_invMixed_0_3[7];
  assign _zz_invMixed_1_37 = (_zz_invMixed_1_19 ^ 8'h1b);
  assign _zz_invMixed_1_38 = 8'h1b;
  assign _zz_invMixed_1_39 = 8'h1b;
  assign _zz_invMixed_2_28 = (_zz_invMixed_2_3[7] ? (_zz_invMixed_2_4 ^ 8'h1b) : _zz_invMixed_2_4);
  assign _zz_invMixed_2_29 = (_zz_invMixed_2_6[7] ? (_zz_invMixed_2_7 ^ 8'h1b) : _zz_invMixed_2_7);
  assign _zz_invMixed_2_30 = _zz_invMixed_2_11[7];
  assign _zz_invMixed_2_31 = (_zz_invMixed_2_12 ^ 8'h1b);
  assign _zz_invMixed_2_32 = _zz_invMixed_2_16[7];
  assign _zz_invMixed_2_33 = (_zz_invMixed_2_17 ^ 8'h1b);
  assign _zz_invMixed_2_34 = _zz_invMixed_2_19[7];
  assign _zz_invMixed_2_35 = (_zz_invMixed_2_20 ^ 8'h1b);
  assign _zz_invMixed_2_36 = 8'h1b;
  assign _zz_invMixed_2_37 = 8'h1b;
  assign _zz_invMixed_2_38 = 8'h1b;
  assign _zz_invMixed_3_28 = (_zz_invMixed_3_3[7] ? (_zz_invMixed_3_4 ^ 8'h1b) : _zz_invMixed_3_4);
  assign _zz_invMixed_3_29 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_3_5 ^ 8'h1b) : _zz_invMixed_3_5);
  assign _zz_invMixed_3_30 = (_zz_invMixed_3_9[7] ? (_zz_invMixed_3_10 ^ 8'h1b) : _zz_invMixed_3_10);
  assign _zz_invMixed_3_31 = (_zz_invMixed_3_12[7] ? (_zz_invMixed_3_13 ^ 8'h1b) : _zz_invMixed_3_13);
  assign _zz_invMixed_3_32 = 8'h1b;
  assign _zz_invMixed_3_33 = 8'h1b;
  assign _zz_invMixed_3_34 = 8'h1b;
  assign _zz_invMixed_4_32 = (_zz_invMixed_4_7[7] ? (_zz_invMixed_4_8 ^ 8'h1b) : _zz_invMixed_4_8);
  assign _zz_invMixed_4_33 = (_zz_invMixed_4_10[7] ? (_zz_invMixed_4_11 ^ 8'h1b) : _zz_invMixed_4_11);
  assign _zz_invMixed_4_34 = _zz_invMixed_4[7];
  assign _zz_invMixed_4_35 = (_zz_invMixed_4_12 ^ 8'h1b);
  assign _zz_invMixed_4_36 = (_zz_invMixed_4_16[7] ? (_zz_invMixed_4_17 ^ 8'h1b) : _zz_invMixed_4_17);
  assign _zz_invMixed_4_37 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_4_18 ^ 8'h1b) : _zz_invMixed_4_18);
  assign _zz_invMixed_4_38 = _zz_invMixed_4_22[7];
  assign _zz_invMixed_4_39 = (_zz_invMixed_4_23 ^ 8'h1b);
  assign _zz_invMixed_4_40 = _zz_invMixed_4_25[7];
  assign _zz_invMixed_4_41 = (_zz_invMixed_4_26 ^ 8'h1b);
  assign _zz_invMixed_5_28 = _zz_invMixed_5_3[7];
  assign _zz_invMixed_5_29 = (_zz_invMixed_5_4 ^ 8'h1b);
  assign _zz_invMixed_5_30 = (_zz_invMixed_5_8[7] ? (_zz_invMixed_5_9 ^ 8'h1b) : _zz_invMixed_5_9);
  assign _zz_invMixed_5_31 = (_zz_invMixed_5_11[7] ? (_zz_invMixed_5_12 ^ 8'h1b) : _zz_invMixed_5_12);
  assign _zz_invMixed_5_32 = _zz_invMixed_4_1[7];
  assign _zz_invMixed_5_33 = (_zz_invMixed_5_13 ^ 8'h1b);
  assign _zz_invMixed_5_34 = _zz_invMixed_5_17[7];
  assign _zz_invMixed_5_35 = (_zz_invMixed_5_18 ^ 8'h1b);
  assign _zz_invMixed_5_36 = _zz_invMixed_4_2[7];
  assign _zz_invMixed_5_37 = (_zz_invMixed_5_19 ^ 8'h1b);
  assign _zz_invMixed_5_38 = 8'h1b;
  assign _zz_invMixed_5_39 = 8'h1b;
  assign _zz_invMixed_6_28 = (_zz_invMixed_6_3[7] ? (_zz_invMixed_6_4 ^ 8'h1b) : _zz_invMixed_6_4);
  assign _zz_invMixed_6_29 = (_zz_invMixed_6_6[7] ? (_zz_invMixed_6_7 ^ 8'h1b) : _zz_invMixed_6_7);
  assign _zz_invMixed_6_30 = _zz_invMixed_6_11[7];
  assign _zz_invMixed_6_31 = (_zz_invMixed_6_12 ^ 8'h1b);
  assign _zz_invMixed_6_32 = _zz_invMixed_6_16[7];
  assign _zz_invMixed_6_33 = (_zz_invMixed_6_17 ^ 8'h1b);
  assign _zz_invMixed_6_34 = _zz_invMixed_6_19[7];
  assign _zz_invMixed_6_35 = (_zz_invMixed_6_20 ^ 8'h1b);
  assign _zz_invMixed_6_36 = 8'h1b;
  assign _zz_invMixed_6_37 = 8'h1b;
  assign _zz_invMixed_6_38 = 8'h1b;
  assign _zz_invMixed_7_28 = (_zz_invMixed_7_3[7] ? (_zz_invMixed_7_4 ^ 8'h1b) : _zz_invMixed_7_4);
  assign _zz_invMixed_7_29 = (_zz_invMixed_4[7] ? (_zz_invMixed_7_5 ^ 8'h1b) : _zz_invMixed_7_5);
  assign _zz_invMixed_7_30 = (_zz_invMixed_7_9[7] ? (_zz_invMixed_7_10 ^ 8'h1b) : _zz_invMixed_7_10);
  assign _zz_invMixed_7_31 = (_zz_invMixed_7_12[7] ? (_zz_invMixed_7_13 ^ 8'h1b) : _zz_invMixed_7_13);
  assign _zz_invMixed_7_32 = 8'h1b;
  assign _zz_invMixed_7_33 = 8'h1b;
  assign _zz_invMixed_7_34 = 8'h1b;
  assign _zz_invMixed_8_32 = (_zz_invMixed_8_7[7] ? (_zz_invMixed_8_8 ^ 8'h1b) : _zz_invMixed_8_8);
  assign _zz_invMixed_8_33 = (_zz_invMixed_8_10[7] ? (_zz_invMixed_8_11 ^ 8'h1b) : _zz_invMixed_8_11);
  assign _zz_invMixed_8_34 = _zz_invMixed_8[7];
  assign _zz_invMixed_8_35 = (_zz_invMixed_8_12 ^ 8'h1b);
  assign _zz_invMixed_8_36 = (_zz_invMixed_8_16[7] ? (_zz_invMixed_8_17 ^ 8'h1b) : _zz_invMixed_8_17);
  assign _zz_invMixed_8_37 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_8_18 ^ 8'h1b) : _zz_invMixed_8_18);
  assign _zz_invMixed_8_38 = _zz_invMixed_8_22[7];
  assign _zz_invMixed_8_39 = (_zz_invMixed_8_23 ^ 8'h1b);
  assign _zz_invMixed_8_40 = _zz_invMixed_8_25[7];
  assign _zz_invMixed_8_41 = (_zz_invMixed_8_26 ^ 8'h1b);
  assign _zz_invMixed_9_28 = _zz_invMixed_9_3[7];
  assign _zz_invMixed_9_29 = (_zz_invMixed_9_4 ^ 8'h1b);
  assign _zz_invMixed_9_30 = (_zz_invMixed_9_8[7] ? (_zz_invMixed_9_9 ^ 8'h1b) : _zz_invMixed_9_9);
  assign _zz_invMixed_9_31 = (_zz_invMixed_9_11[7] ? (_zz_invMixed_9_12 ^ 8'h1b) : _zz_invMixed_9_12);
  assign _zz_invMixed_9_32 = _zz_invMixed_8_1[7];
  assign _zz_invMixed_9_33 = (_zz_invMixed_9_13 ^ 8'h1b);
  assign _zz_invMixed_9_34 = _zz_invMixed_9_17[7];
  assign _zz_invMixed_9_35 = (_zz_invMixed_9_18 ^ 8'h1b);
  assign _zz_invMixed_9_36 = _zz_invMixed_8_2[7];
  assign _zz_invMixed_9_37 = (_zz_invMixed_9_19 ^ 8'h1b);
  assign _zz_invMixed_9_38 = 8'h1b;
  assign _zz_invMixed_9_39 = 8'h1b;
  assign _zz_invMixed_10_28 = (_zz_invMixed_10_3[7] ? (_zz_invMixed_10_4 ^ 8'h1b) : _zz_invMixed_10_4);
  assign _zz_invMixed_10_29 = (_zz_invMixed_10_6[7] ? (_zz_invMixed_10_7 ^ 8'h1b) : _zz_invMixed_10_7);
  assign _zz_invMixed_10_30 = _zz_invMixed_10_11[7];
  assign _zz_invMixed_10_31 = (_zz_invMixed_10_12 ^ 8'h1b);
  assign _zz_invMixed_10_32 = _zz_invMixed_10_16[7];
  assign _zz_invMixed_10_33 = (_zz_invMixed_10_17 ^ 8'h1b);
  assign _zz_invMixed_10_34 = _zz_invMixed_10_19[7];
  assign _zz_invMixed_10_35 = (_zz_invMixed_10_20 ^ 8'h1b);
  assign _zz_invMixed_10_36 = 8'h1b;
  assign _zz_invMixed_10_37 = 8'h1b;
  assign _zz_invMixed_10_38 = 8'h1b;
  assign _zz_invMixed_11_28 = (_zz_invMixed_11_3[7] ? (_zz_invMixed_11_4 ^ 8'h1b) : _zz_invMixed_11_4);
  assign _zz_invMixed_11_29 = (_zz_invMixed_8[7] ? (_zz_invMixed_11_5 ^ 8'h1b) : _zz_invMixed_11_5);
  assign _zz_invMixed_11_30 = (_zz_invMixed_11_9[7] ? (_zz_invMixed_11_10 ^ 8'h1b) : _zz_invMixed_11_10);
  assign _zz_invMixed_11_31 = (_zz_invMixed_11_12[7] ? (_zz_invMixed_11_13 ^ 8'h1b) : _zz_invMixed_11_13);
  assign _zz_invMixed_11_32 = 8'h1b;
  assign _zz_invMixed_11_33 = 8'h1b;
  assign _zz_invMixed_11_34 = 8'h1b;
  assign _zz_invMixed_12_32 = (_zz_invMixed_12_7[7] ? (_zz_invMixed_12_8 ^ 8'h1b) : _zz_invMixed_12_8);
  assign _zz_invMixed_12_33 = (_zz_invMixed_12_10[7] ? (_zz_invMixed_12_11 ^ 8'h1b) : _zz_invMixed_12_11);
  assign _zz_invMixed_12_34 = _zz_invMixed_12[7];
  assign _zz_invMixed_12_35 = (_zz_invMixed_12_12 ^ 8'h1b);
  assign _zz_invMixed_12_36 = (_zz_invMixed_12_16[7] ? (_zz_invMixed_12_17 ^ 8'h1b) : _zz_invMixed_12_17);
  assign _zz_invMixed_12_37 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_12_18 ^ 8'h1b) : _zz_invMixed_12_18);
  assign _zz_invMixed_12_38 = _zz_invMixed_12_22[7];
  assign _zz_invMixed_12_39 = (_zz_invMixed_12_23 ^ 8'h1b);
  assign _zz_invMixed_12_40 = _zz_invMixed_12_25[7];
  assign _zz_invMixed_12_41 = (_zz_invMixed_12_26 ^ 8'h1b);
  assign _zz_invMixed_13_28 = _zz_invMixed_13_3[7];
  assign _zz_invMixed_13_29 = (_zz_invMixed_13_4 ^ 8'h1b);
  assign _zz_invMixed_13_30 = (_zz_invMixed_13_8[7] ? (_zz_invMixed_13_9 ^ 8'h1b) : _zz_invMixed_13_9);
  assign _zz_invMixed_13_31 = (_zz_invMixed_13_11[7] ? (_zz_invMixed_13_12 ^ 8'h1b) : _zz_invMixed_13_12);
  assign _zz_invMixed_13_32 = _zz_invMixed_12_1[7];
  assign _zz_invMixed_13_33 = (_zz_invMixed_13_13 ^ 8'h1b);
  assign _zz_invMixed_13_34 = _zz_invMixed_13_17[7];
  assign _zz_invMixed_13_35 = (_zz_invMixed_13_18 ^ 8'h1b);
  assign _zz_invMixed_13_36 = _zz_invMixed_12_2[7];
  assign _zz_invMixed_13_37 = (_zz_invMixed_13_19 ^ 8'h1b);
  assign _zz_invMixed_13_38 = 8'h1b;
  assign _zz_invMixed_13_39 = 8'h1b;
  assign _zz_invMixed_14_28 = (_zz_invMixed_14_3[7] ? (_zz_invMixed_14_4 ^ 8'h1b) : _zz_invMixed_14_4);
  assign _zz_invMixed_14_29 = (_zz_invMixed_14_6[7] ? (_zz_invMixed_14_7 ^ 8'h1b) : _zz_invMixed_14_7);
  assign _zz_invMixed_14_30 = _zz_invMixed_14_11[7];
  assign _zz_invMixed_14_31 = (_zz_invMixed_14_12 ^ 8'h1b);
  assign _zz_invMixed_14_32 = _zz_invMixed_14_16[7];
  assign _zz_invMixed_14_33 = (_zz_invMixed_14_17 ^ 8'h1b);
  assign _zz_invMixed_14_34 = _zz_invMixed_14_19[7];
  assign _zz_invMixed_14_35 = (_zz_invMixed_14_20 ^ 8'h1b);
  assign _zz_invMixed_14_36 = 8'h1b;
  assign _zz_invMixed_14_37 = 8'h1b;
  assign _zz_invMixed_14_38 = 8'h1b;
  assign _zz_invMixed_15_28 = (_zz_invMixed_15_3[7] ? (_zz_invMixed_15_4 ^ 8'h1b) : _zz_invMixed_15_4);
  assign _zz_invMixed_15_29 = (_zz_invMixed_12[7] ? (_zz_invMixed_15_5 ^ 8'h1b) : _zz_invMixed_15_5);
  assign _zz_invMixed_15_30 = (_zz_invMixed_15_9[7] ? (_zz_invMixed_15_10 ^ 8'h1b) : _zz_invMixed_15_10);
  assign _zz_invMixed_15_31 = (_zz_invMixed_15_12[7] ? (_zz_invMixed_15_13 ^ 8'h1b) : _zz_invMixed_15_13);
  assign _zz_invMixed_15_32 = 8'h1b;
  assign _zz_invMixed_15_33 = 8'h1b;
  assign _zz_invMixed_15_34 = 8'h1b;
  assign _zz_stateReg_95 = {{{{invMixed_0,invMixed_1},invMixed_2},invMixed_3},invMixed_4};
  assign _zz_stateReg_96 = invMixed_5;
  always @(*) begin
    case(_zz__zz_stateReg_4_1)
      8'b00000000 : _zz__zz_stateReg_4 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_4 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_4 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_4 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_4 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_4 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_4 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_4 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_4 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_4 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_4 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_4 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_4 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_4 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_4 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_4 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_4 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_4 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_4 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_4 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_4 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_4 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_4 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_4 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_4 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_4 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_4 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_4 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_4 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_4 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_4 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_4 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_4 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_4 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_4 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_4 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_4 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_4 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_4 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_4 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_4 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_4 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_4 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_4 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_4 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_4 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_4 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_4 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_4 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_4 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_4 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_4 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_4 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_4 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_4 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_4 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_4 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_4 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_4 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_4 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_4 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_4 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_4 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_4 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_4 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_4 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_4 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_4 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_4 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_4 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_4 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_4 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_4 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_4 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_4 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_4 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_4 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_4 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_4 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_4 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_4 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_4 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_4 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_4 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_4 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_4 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_4 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_4 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_4 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_4 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_4 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_4 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_4 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_4 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_4 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_4 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_4 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_4 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_4 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_4 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_4 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_4 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_4 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_4 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_4 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_4 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_4 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_4 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_4 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_4 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_4 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_4 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_4 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_4 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_4 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_4 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_4 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_4 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_4 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_4 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_4 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_4 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_4 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_4 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_4 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_4 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_4 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_4 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_4 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_4 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_4 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_4 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_4 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_4 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_4 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_4 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_4 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_4 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_4 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_4 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_4 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_4 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_4 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_4 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_4 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_4 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_4 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_4 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_4 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_4 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_4 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_4 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_4 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_4 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_4 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_4 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_4 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_4 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_4 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_4 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_4 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_4 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_4 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_4 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_4 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_4 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_4 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_4 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_4 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_4 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_4 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_4 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_4 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_4 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_4 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_4 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_4 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_4 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_4 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_4 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_4 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_4 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_4 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_4 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_4 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_4 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_4 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_4 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_4 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_4 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_4 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_4 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_4 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_4 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_4 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_4 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_4 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_4 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_4 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_4 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_4 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_4 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_4 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_4 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_4 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_4 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_4 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_4 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_4 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_4 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_4 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_4 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_4 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_4 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_4 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_4 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_4 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_4 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_4 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_4 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_4 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_4 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_4 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_4 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_4 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_4 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_4 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_4 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_4 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_4 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_4 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_4 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_4 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_4 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_4 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_4 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_4 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_4 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_4 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_4 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_4 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_4 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_4 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_4 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_4 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_4 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_4 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_4 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_4 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_4 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_4 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_4 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_4 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_4 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_4 = sboxRom_254;
      default : _zz__zz_stateReg_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_8_1)
      8'b00000000 : _zz__zz_stateReg_8 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_8 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_8 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_8 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_8 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_8 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_8 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_8 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_8 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_8 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_8 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_8 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_8 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_8 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_8 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_8 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_8 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_8 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_8 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_8 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_8 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_8 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_8 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_8 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_8 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_8 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_8 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_8 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_8 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_8 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_8 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_8 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_8 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_8 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_8 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_8 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_8 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_8 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_8 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_8 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_8 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_8 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_8 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_8 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_8 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_8 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_8 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_8 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_8 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_8 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_8 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_8 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_8 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_8 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_8 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_8 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_8 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_8 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_8 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_8 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_8 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_8 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_8 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_8 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_8 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_8 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_8 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_8 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_8 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_8 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_8 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_8 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_8 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_8 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_8 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_8 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_8 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_8 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_8 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_8 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_8 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_8 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_8 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_8 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_8 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_8 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_8 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_8 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_8 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_8 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_8 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_8 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_8 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_8 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_8 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_8 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_8 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_8 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_8 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_8 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_8 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_8 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_8 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_8 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_8 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_8 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_8 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_8 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_8 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_8 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_8 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_8 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_8 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_8 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_8 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_8 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_8 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_8 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_8 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_8 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_8 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_8 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_8 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_8 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_8 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_8 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_8 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_8 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_8 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_8 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_8 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_8 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_8 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_8 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_8 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_8 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_8 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_8 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_8 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_8 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_8 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_8 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_8 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_8 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_8 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_8 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_8 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_8 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_8 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_8 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_8 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_8 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_8 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_8 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_8 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_8 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_8 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_8 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_8 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_8 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_8 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_8 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_8 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_8 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_8 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_8 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_8 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_8 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_8 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_8 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_8 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_8 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_8 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_8 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_8 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_8 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_8 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_8 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_8 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_8 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_8 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_8 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_8 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_8 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_8 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_8 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_8 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_8 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_8 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_8 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_8 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_8 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_8 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_8 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_8 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_8 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_8 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_8 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_8 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_8 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_8 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_8 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_8 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_8 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_8 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_8 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_8 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_8 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_8 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_8 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_8 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_8 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_8 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_8 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_8 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_8 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_8 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_8 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_8 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_8 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_8 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_8 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_8 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_8 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_8 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_8 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_8 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_8 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_8 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_8 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_8 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_8 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_8 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_8 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_8 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_8 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_8 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_8 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_8 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_8 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_8 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_8 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_8 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_8 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_8 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_8 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_8 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_8 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_8 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_8 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_8 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_8 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_8 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_8 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_8 = sboxRom_254;
      default : _zz__zz_stateReg_8 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_12_1)
      8'b00000000 : _zz__zz_stateReg_12 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_12 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_12 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_12 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_12 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_12 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_12 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_12 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_12 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_12 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_12 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_12 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_12 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_12 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_12 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_12 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_12 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_12 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_12 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_12 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_12 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_12 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_12 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_12 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_12 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_12 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_12 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_12 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_12 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_12 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_12 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_12 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_12 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_12 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_12 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_12 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_12 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_12 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_12 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_12 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_12 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_12 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_12 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_12 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_12 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_12 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_12 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_12 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_12 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_12 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_12 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_12 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_12 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_12 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_12 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_12 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_12 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_12 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_12 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_12 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_12 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_12 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_12 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_12 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_12 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_12 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_12 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_12 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_12 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_12 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_12 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_12 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_12 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_12 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_12 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_12 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_12 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_12 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_12 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_12 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_12 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_12 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_12 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_12 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_12 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_12 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_12 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_12 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_12 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_12 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_12 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_12 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_12 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_12 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_12 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_12 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_12 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_12 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_12 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_12 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_12 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_12 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_12 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_12 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_12 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_12 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_12 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_12 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_12 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_12 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_12 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_12 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_12 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_12 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_12 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_12 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_12 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_12 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_12 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_12 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_12 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_12 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_12 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_12 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_12 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_12 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_12 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_12 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_12 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_12 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_12 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_12 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_12 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_12 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_12 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_12 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_12 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_12 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_12 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_12 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_12 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_12 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_12 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_12 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_12 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_12 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_12 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_12 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_12 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_12 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_12 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_12 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_12 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_12 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_12 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_12 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_12 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_12 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_12 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_12 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_12 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_12 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_12 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_12 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_12 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_12 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_12 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_12 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_12 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_12 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_12 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_12 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_12 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_12 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_12 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_12 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_12 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_12 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_12 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_12 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_12 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_12 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_12 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_12 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_12 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_12 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_12 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_12 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_12 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_12 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_12 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_12 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_12 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_12 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_12 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_12 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_12 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_12 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_12 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_12 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_12 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_12 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_12 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_12 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_12 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_12 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_12 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_12 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_12 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_12 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_12 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_12 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_12 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_12 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_12 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_12 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_12 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_12 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_12 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_12 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_12 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_12 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_12 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_12 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_12 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_12 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_12 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_12 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_12 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_12 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_12 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_12 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_12 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_12 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_12 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_12 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_12 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_12 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_12 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_12 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_12 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_12 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_12 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_12 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_12 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_12 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_12 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_12 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_12 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_12 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_12 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_12 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_12 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_12 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_12 = sboxRom_254;
      default : _zz__zz_stateReg_12 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_16_1)
      8'b00000000 : _zz__zz_stateReg_16 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_16 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_16 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_16 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_16 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_16 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_16 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_16 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_16 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_16 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_16 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_16 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_16 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_16 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_16 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_16 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_16 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_16 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_16 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_16 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_16 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_16 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_16 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_16 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_16 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_16 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_16 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_16 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_16 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_16 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_16 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_16 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_16 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_16 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_16 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_16 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_16 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_16 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_16 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_16 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_16 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_16 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_16 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_16 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_16 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_16 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_16 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_16 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_16 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_16 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_16 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_16 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_16 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_16 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_16 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_16 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_16 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_16 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_16 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_16 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_16 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_16 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_16 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_16 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_16 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_16 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_16 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_16 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_16 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_16 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_16 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_16 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_16 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_16 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_16 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_16 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_16 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_16 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_16 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_16 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_16 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_16 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_16 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_16 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_16 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_16 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_16 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_16 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_16 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_16 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_16 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_16 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_16 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_16 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_16 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_16 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_16 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_16 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_16 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_16 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_16 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_16 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_16 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_16 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_16 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_16 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_16 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_16 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_16 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_16 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_16 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_16 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_16 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_16 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_16 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_16 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_16 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_16 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_16 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_16 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_16 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_16 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_16 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_16 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_16 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_16 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_16 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_16 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_16 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_16 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_16 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_16 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_16 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_16 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_16 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_16 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_16 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_16 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_16 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_16 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_16 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_16 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_16 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_16 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_16 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_16 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_16 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_16 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_16 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_16 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_16 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_16 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_16 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_16 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_16 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_16 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_16 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_16 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_16 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_16 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_16 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_16 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_16 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_16 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_16 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_16 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_16 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_16 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_16 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_16 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_16 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_16 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_16 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_16 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_16 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_16 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_16 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_16 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_16 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_16 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_16 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_16 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_16 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_16 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_16 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_16 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_16 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_16 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_16 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_16 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_16 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_16 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_16 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_16 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_16 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_16 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_16 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_16 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_16 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_16 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_16 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_16 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_16 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_16 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_16 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_16 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_16 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_16 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_16 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_16 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_16 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_16 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_16 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_16 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_16 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_16 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_16 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_16 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_16 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_16 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_16 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_16 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_16 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_16 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_16 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_16 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_16 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_16 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_16 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_16 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_16 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_16 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_16 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_16 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_16 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_16 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_16 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_16 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_16 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_16 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_16 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_16 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_16 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_16 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_16 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_16 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_16 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_16 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_16 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_16 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_16 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_16 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_16 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_16 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_16 = sboxRom_254;
      default : _zz__zz_stateReg_16 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_5_1)
      8'b00000000 : _zz__zz_stateReg_5 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_5 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_5 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_5 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_5 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_5 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_5 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_5 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_5 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_5 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_5 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_5 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_5 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_5 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_5 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_5 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_5 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_5 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_5 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_5 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_5 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_5 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_5 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_5 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_5 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_5 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_5 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_5 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_5 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_5 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_5 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_5 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_5 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_5 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_5 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_5 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_5 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_5 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_5 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_5 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_5 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_5 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_5 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_5 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_5 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_5 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_5 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_5 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_5 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_5 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_5 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_5 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_5 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_5 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_5 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_5 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_5 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_5 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_5 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_5 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_5 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_5 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_5 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_5 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_5 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_5 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_5 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_5 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_5 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_5 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_5 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_5 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_5 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_5 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_5 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_5 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_5 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_5 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_5 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_5 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_5 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_5 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_5 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_5 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_5 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_5 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_5 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_5 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_5 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_5 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_5 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_5 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_5 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_5 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_5 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_5 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_5 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_5 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_5 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_5 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_5 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_5 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_5 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_5 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_5 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_5 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_5 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_5 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_5 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_5 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_5 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_5 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_5 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_5 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_5 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_5 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_5 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_5 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_5 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_5 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_5 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_5 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_5 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_5 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_5 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_5 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_5 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_5 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_5 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_5 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_5 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_5 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_5 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_5 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_5 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_5 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_5 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_5 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_5 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_5 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_5 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_5 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_5 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_5 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_5 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_5 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_5 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_5 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_5 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_5 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_5 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_5 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_5 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_5 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_5 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_5 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_5 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_5 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_5 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_5 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_5 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_5 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_5 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_5 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_5 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_5 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_5 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_5 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_5 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_5 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_5 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_5 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_5 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_5 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_5 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_5 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_5 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_5 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_5 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_5 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_5 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_5 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_5 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_5 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_5 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_5 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_5 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_5 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_5 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_5 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_5 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_5 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_5 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_5 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_5 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_5 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_5 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_5 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_5 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_5 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_5 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_5 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_5 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_5 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_5 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_5 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_5 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_5 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_5 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_5 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_5 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_5 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_5 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_5 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_5 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_5 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_5 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_5 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_5 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_5 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_5 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_5 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_5 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_5 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_5 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_5 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_5 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_5 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_5 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_5 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_5 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_5 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_5 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_5 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_5 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_5 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_5 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_5 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_5 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_5 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_5 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_5 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_5 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_5 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_5 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_5 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_5 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_5 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_5 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_5 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_5 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_5 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_5 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_5 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_5 = sboxRom_254;
      default : _zz__zz_stateReg_5 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_9_1)
      8'b00000000 : _zz__zz_stateReg_9 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_9 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_9 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_9 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_9 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_9 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_9 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_9 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_9 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_9 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_9 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_9 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_9 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_9 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_9 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_9 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_9 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_9 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_9 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_9 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_9 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_9 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_9 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_9 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_9 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_9 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_9 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_9 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_9 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_9 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_9 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_9 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_9 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_9 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_9 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_9 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_9 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_9 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_9 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_9 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_9 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_9 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_9 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_9 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_9 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_9 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_9 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_9 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_9 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_9 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_9 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_9 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_9 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_9 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_9 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_9 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_9 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_9 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_9 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_9 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_9 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_9 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_9 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_9 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_9 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_9 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_9 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_9 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_9 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_9 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_9 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_9 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_9 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_9 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_9 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_9 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_9 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_9 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_9 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_9 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_9 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_9 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_9 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_9 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_9 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_9 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_9 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_9 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_9 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_9 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_9 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_9 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_9 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_9 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_9 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_9 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_9 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_9 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_9 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_9 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_9 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_9 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_9 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_9 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_9 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_9 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_9 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_9 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_9 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_9 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_9 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_9 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_9 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_9 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_9 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_9 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_9 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_9 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_9 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_9 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_9 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_9 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_9 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_9 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_9 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_9 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_9 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_9 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_9 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_9 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_9 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_9 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_9 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_9 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_9 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_9 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_9 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_9 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_9 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_9 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_9 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_9 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_9 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_9 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_9 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_9 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_9 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_9 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_9 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_9 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_9 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_9 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_9 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_9 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_9 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_9 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_9 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_9 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_9 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_9 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_9 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_9 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_9 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_9 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_9 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_9 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_9 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_9 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_9 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_9 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_9 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_9 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_9 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_9 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_9 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_9 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_9 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_9 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_9 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_9 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_9 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_9 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_9 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_9 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_9 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_9 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_9 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_9 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_9 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_9 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_9 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_9 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_9 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_9 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_9 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_9 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_9 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_9 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_9 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_9 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_9 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_9 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_9 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_9 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_9 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_9 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_9 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_9 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_9 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_9 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_9 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_9 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_9 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_9 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_9 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_9 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_9 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_9 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_9 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_9 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_9 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_9 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_9 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_9 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_9 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_9 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_9 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_9 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_9 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_9 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_9 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_9 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_9 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_9 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_9 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_9 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_9 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_9 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_9 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_9 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_9 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_9 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_9 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_9 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_9 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_9 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_9 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_9 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_9 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_9 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_9 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_9 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_9 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_9 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_9 = sboxRom_254;
      default : _zz__zz_stateReg_9 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_13_1)
      8'b00000000 : _zz__zz_stateReg_13 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_13 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_13 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_13 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_13 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_13 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_13 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_13 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_13 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_13 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_13 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_13 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_13 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_13 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_13 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_13 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_13 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_13 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_13 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_13 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_13 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_13 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_13 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_13 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_13 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_13 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_13 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_13 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_13 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_13 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_13 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_13 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_13 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_13 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_13 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_13 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_13 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_13 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_13 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_13 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_13 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_13 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_13 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_13 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_13 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_13 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_13 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_13 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_13 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_13 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_13 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_13 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_13 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_13 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_13 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_13 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_13 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_13 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_13 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_13 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_13 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_13 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_13 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_13 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_13 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_13 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_13 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_13 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_13 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_13 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_13 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_13 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_13 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_13 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_13 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_13 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_13 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_13 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_13 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_13 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_13 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_13 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_13 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_13 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_13 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_13 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_13 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_13 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_13 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_13 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_13 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_13 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_13 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_13 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_13 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_13 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_13 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_13 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_13 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_13 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_13 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_13 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_13 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_13 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_13 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_13 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_13 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_13 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_13 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_13 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_13 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_13 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_13 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_13 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_13 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_13 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_13 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_13 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_13 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_13 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_13 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_13 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_13 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_13 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_13 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_13 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_13 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_13 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_13 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_13 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_13 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_13 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_13 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_13 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_13 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_13 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_13 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_13 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_13 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_13 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_13 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_13 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_13 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_13 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_13 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_13 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_13 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_13 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_13 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_13 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_13 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_13 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_13 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_13 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_13 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_13 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_13 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_13 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_13 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_13 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_13 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_13 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_13 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_13 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_13 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_13 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_13 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_13 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_13 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_13 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_13 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_13 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_13 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_13 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_13 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_13 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_13 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_13 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_13 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_13 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_13 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_13 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_13 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_13 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_13 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_13 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_13 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_13 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_13 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_13 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_13 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_13 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_13 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_13 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_13 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_13 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_13 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_13 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_13 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_13 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_13 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_13 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_13 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_13 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_13 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_13 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_13 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_13 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_13 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_13 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_13 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_13 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_13 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_13 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_13 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_13 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_13 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_13 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_13 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_13 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_13 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_13 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_13 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_13 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_13 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_13 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_13 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_13 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_13 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_13 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_13 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_13 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_13 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_13 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_13 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_13 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_13 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_13 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_13 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_13 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_13 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_13 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_13 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_13 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_13 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_13 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_13 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_13 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_13 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_13 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_13 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_13 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_13 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_13 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_13 = sboxRom_254;
      default : _zz__zz_stateReg_13 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_17_1)
      8'b00000000 : _zz__zz_stateReg_17 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_17 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_17 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_17 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_17 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_17 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_17 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_17 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_17 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_17 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_17 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_17 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_17 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_17 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_17 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_17 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_17 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_17 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_17 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_17 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_17 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_17 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_17 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_17 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_17 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_17 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_17 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_17 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_17 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_17 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_17 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_17 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_17 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_17 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_17 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_17 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_17 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_17 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_17 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_17 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_17 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_17 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_17 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_17 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_17 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_17 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_17 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_17 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_17 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_17 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_17 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_17 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_17 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_17 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_17 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_17 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_17 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_17 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_17 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_17 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_17 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_17 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_17 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_17 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_17 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_17 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_17 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_17 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_17 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_17 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_17 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_17 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_17 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_17 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_17 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_17 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_17 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_17 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_17 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_17 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_17 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_17 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_17 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_17 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_17 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_17 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_17 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_17 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_17 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_17 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_17 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_17 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_17 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_17 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_17 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_17 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_17 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_17 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_17 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_17 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_17 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_17 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_17 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_17 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_17 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_17 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_17 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_17 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_17 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_17 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_17 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_17 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_17 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_17 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_17 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_17 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_17 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_17 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_17 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_17 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_17 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_17 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_17 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_17 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_17 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_17 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_17 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_17 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_17 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_17 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_17 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_17 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_17 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_17 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_17 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_17 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_17 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_17 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_17 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_17 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_17 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_17 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_17 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_17 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_17 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_17 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_17 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_17 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_17 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_17 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_17 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_17 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_17 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_17 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_17 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_17 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_17 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_17 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_17 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_17 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_17 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_17 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_17 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_17 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_17 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_17 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_17 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_17 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_17 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_17 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_17 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_17 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_17 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_17 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_17 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_17 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_17 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_17 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_17 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_17 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_17 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_17 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_17 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_17 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_17 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_17 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_17 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_17 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_17 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_17 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_17 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_17 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_17 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_17 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_17 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_17 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_17 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_17 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_17 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_17 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_17 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_17 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_17 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_17 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_17 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_17 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_17 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_17 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_17 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_17 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_17 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_17 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_17 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_17 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_17 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_17 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_17 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_17 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_17 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_17 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_17 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_17 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_17 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_17 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_17 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_17 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_17 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_17 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_17 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_17 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_17 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_17 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_17 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_17 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_17 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_17 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_17 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_17 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_17 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_17 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_17 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_17 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_17 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_17 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_17 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_17 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_17 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_17 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_17 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_17 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_17 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_17 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_17 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_17 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_17 = sboxRom_254;
      default : _zz__zz_stateReg_17 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_6_1)
      8'b00000000 : _zz__zz_stateReg_6 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_6 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_6 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_6 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_6 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_6 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_6 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_6 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_6 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_6 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_6 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_6 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_6 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_6 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_6 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_6 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_6 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_6 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_6 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_6 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_6 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_6 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_6 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_6 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_6 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_6 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_6 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_6 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_6 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_6 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_6 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_6 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_6 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_6 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_6 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_6 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_6 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_6 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_6 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_6 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_6 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_6 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_6 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_6 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_6 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_6 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_6 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_6 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_6 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_6 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_6 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_6 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_6 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_6 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_6 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_6 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_6 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_6 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_6 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_6 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_6 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_6 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_6 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_6 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_6 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_6 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_6 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_6 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_6 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_6 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_6 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_6 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_6 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_6 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_6 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_6 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_6 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_6 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_6 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_6 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_6 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_6 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_6 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_6 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_6 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_6 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_6 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_6 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_6 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_6 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_6 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_6 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_6 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_6 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_6 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_6 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_6 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_6 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_6 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_6 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_6 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_6 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_6 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_6 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_6 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_6 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_6 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_6 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_6 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_6 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_6 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_6 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_6 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_6 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_6 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_6 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_6 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_6 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_6 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_6 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_6 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_6 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_6 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_6 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_6 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_6 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_6 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_6 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_6 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_6 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_6 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_6 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_6 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_6 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_6 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_6 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_6 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_6 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_6 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_6 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_6 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_6 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_6 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_6 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_6 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_6 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_6 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_6 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_6 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_6 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_6 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_6 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_6 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_6 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_6 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_6 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_6 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_6 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_6 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_6 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_6 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_6 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_6 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_6 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_6 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_6 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_6 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_6 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_6 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_6 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_6 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_6 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_6 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_6 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_6 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_6 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_6 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_6 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_6 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_6 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_6 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_6 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_6 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_6 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_6 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_6 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_6 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_6 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_6 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_6 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_6 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_6 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_6 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_6 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_6 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_6 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_6 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_6 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_6 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_6 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_6 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_6 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_6 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_6 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_6 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_6 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_6 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_6 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_6 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_6 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_6 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_6 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_6 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_6 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_6 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_6 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_6 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_6 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_6 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_6 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_6 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_6 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_6 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_6 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_6 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_6 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_6 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_6 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_6 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_6 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_6 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_6 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_6 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_6 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_6 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_6 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_6 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_6 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_6 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_6 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_6 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_6 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_6 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_6 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_6 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_6 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_6 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_6 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_6 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_6 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_6 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_6 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_6 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_6 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_6 = sboxRom_254;
      default : _zz__zz_stateReg_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_10_1)
      8'b00000000 : _zz__zz_stateReg_10 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_10 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_10 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_10 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_10 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_10 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_10 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_10 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_10 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_10 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_10 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_10 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_10 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_10 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_10 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_10 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_10 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_10 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_10 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_10 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_10 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_10 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_10 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_10 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_10 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_10 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_10 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_10 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_10 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_10 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_10 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_10 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_10 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_10 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_10 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_10 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_10 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_10 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_10 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_10 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_10 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_10 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_10 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_10 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_10 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_10 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_10 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_10 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_10 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_10 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_10 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_10 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_10 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_10 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_10 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_10 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_10 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_10 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_10 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_10 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_10 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_10 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_10 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_10 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_10 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_10 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_10 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_10 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_10 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_10 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_10 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_10 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_10 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_10 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_10 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_10 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_10 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_10 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_10 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_10 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_10 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_10 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_10 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_10 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_10 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_10 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_10 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_10 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_10 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_10 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_10 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_10 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_10 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_10 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_10 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_10 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_10 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_10 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_10 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_10 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_10 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_10 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_10 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_10 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_10 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_10 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_10 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_10 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_10 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_10 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_10 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_10 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_10 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_10 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_10 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_10 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_10 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_10 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_10 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_10 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_10 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_10 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_10 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_10 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_10 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_10 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_10 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_10 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_10 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_10 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_10 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_10 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_10 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_10 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_10 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_10 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_10 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_10 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_10 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_10 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_10 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_10 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_10 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_10 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_10 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_10 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_10 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_10 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_10 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_10 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_10 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_10 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_10 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_10 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_10 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_10 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_10 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_10 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_10 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_10 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_10 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_10 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_10 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_10 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_10 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_10 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_10 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_10 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_10 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_10 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_10 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_10 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_10 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_10 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_10 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_10 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_10 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_10 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_10 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_10 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_10 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_10 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_10 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_10 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_10 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_10 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_10 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_10 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_10 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_10 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_10 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_10 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_10 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_10 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_10 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_10 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_10 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_10 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_10 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_10 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_10 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_10 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_10 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_10 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_10 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_10 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_10 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_10 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_10 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_10 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_10 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_10 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_10 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_10 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_10 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_10 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_10 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_10 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_10 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_10 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_10 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_10 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_10 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_10 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_10 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_10 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_10 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_10 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_10 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_10 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_10 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_10 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_10 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_10 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_10 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_10 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_10 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_10 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_10 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_10 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_10 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_10 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_10 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_10 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_10 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_10 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_10 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_10 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_10 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_10 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_10 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_10 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_10 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_10 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_10 = sboxRom_254;
      default : _zz__zz_stateReg_10 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_14_1)
      8'b00000000 : _zz__zz_stateReg_14 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_14 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_14 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_14 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_14 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_14 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_14 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_14 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_14 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_14 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_14 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_14 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_14 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_14 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_14 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_14 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_14 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_14 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_14 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_14 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_14 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_14 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_14 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_14 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_14 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_14 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_14 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_14 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_14 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_14 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_14 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_14 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_14 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_14 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_14 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_14 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_14 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_14 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_14 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_14 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_14 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_14 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_14 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_14 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_14 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_14 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_14 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_14 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_14 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_14 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_14 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_14 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_14 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_14 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_14 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_14 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_14 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_14 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_14 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_14 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_14 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_14 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_14 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_14 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_14 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_14 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_14 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_14 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_14 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_14 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_14 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_14 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_14 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_14 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_14 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_14 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_14 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_14 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_14 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_14 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_14 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_14 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_14 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_14 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_14 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_14 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_14 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_14 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_14 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_14 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_14 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_14 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_14 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_14 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_14 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_14 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_14 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_14 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_14 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_14 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_14 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_14 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_14 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_14 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_14 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_14 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_14 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_14 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_14 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_14 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_14 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_14 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_14 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_14 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_14 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_14 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_14 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_14 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_14 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_14 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_14 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_14 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_14 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_14 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_14 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_14 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_14 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_14 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_14 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_14 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_14 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_14 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_14 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_14 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_14 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_14 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_14 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_14 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_14 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_14 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_14 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_14 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_14 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_14 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_14 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_14 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_14 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_14 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_14 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_14 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_14 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_14 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_14 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_14 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_14 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_14 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_14 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_14 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_14 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_14 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_14 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_14 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_14 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_14 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_14 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_14 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_14 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_14 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_14 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_14 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_14 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_14 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_14 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_14 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_14 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_14 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_14 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_14 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_14 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_14 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_14 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_14 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_14 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_14 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_14 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_14 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_14 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_14 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_14 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_14 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_14 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_14 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_14 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_14 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_14 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_14 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_14 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_14 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_14 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_14 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_14 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_14 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_14 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_14 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_14 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_14 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_14 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_14 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_14 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_14 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_14 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_14 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_14 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_14 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_14 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_14 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_14 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_14 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_14 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_14 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_14 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_14 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_14 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_14 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_14 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_14 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_14 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_14 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_14 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_14 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_14 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_14 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_14 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_14 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_14 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_14 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_14 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_14 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_14 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_14 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_14 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_14 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_14 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_14 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_14 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_14 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_14 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_14 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_14 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_14 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_14 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_14 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_14 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_14 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_14 = sboxRom_254;
      default : _zz__zz_stateReg_14 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_18_1)
      8'b00000000 : _zz__zz_stateReg_18 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_18 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_18 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_18 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_18 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_18 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_18 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_18 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_18 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_18 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_18 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_18 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_18 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_18 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_18 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_18 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_18 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_18 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_18 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_18 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_18 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_18 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_18 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_18 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_18 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_18 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_18 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_18 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_18 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_18 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_18 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_18 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_18 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_18 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_18 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_18 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_18 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_18 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_18 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_18 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_18 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_18 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_18 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_18 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_18 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_18 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_18 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_18 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_18 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_18 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_18 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_18 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_18 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_18 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_18 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_18 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_18 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_18 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_18 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_18 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_18 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_18 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_18 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_18 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_18 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_18 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_18 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_18 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_18 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_18 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_18 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_18 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_18 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_18 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_18 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_18 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_18 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_18 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_18 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_18 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_18 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_18 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_18 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_18 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_18 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_18 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_18 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_18 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_18 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_18 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_18 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_18 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_18 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_18 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_18 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_18 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_18 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_18 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_18 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_18 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_18 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_18 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_18 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_18 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_18 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_18 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_18 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_18 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_18 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_18 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_18 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_18 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_18 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_18 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_18 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_18 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_18 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_18 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_18 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_18 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_18 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_18 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_18 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_18 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_18 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_18 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_18 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_18 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_18 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_18 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_18 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_18 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_18 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_18 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_18 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_18 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_18 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_18 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_18 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_18 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_18 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_18 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_18 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_18 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_18 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_18 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_18 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_18 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_18 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_18 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_18 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_18 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_18 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_18 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_18 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_18 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_18 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_18 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_18 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_18 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_18 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_18 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_18 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_18 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_18 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_18 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_18 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_18 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_18 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_18 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_18 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_18 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_18 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_18 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_18 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_18 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_18 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_18 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_18 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_18 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_18 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_18 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_18 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_18 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_18 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_18 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_18 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_18 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_18 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_18 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_18 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_18 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_18 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_18 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_18 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_18 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_18 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_18 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_18 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_18 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_18 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_18 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_18 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_18 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_18 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_18 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_18 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_18 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_18 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_18 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_18 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_18 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_18 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_18 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_18 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_18 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_18 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_18 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_18 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_18 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_18 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_18 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_18 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_18 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_18 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_18 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_18 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_18 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_18 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_18 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_18 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_18 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_18 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_18 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_18 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_18 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_18 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_18 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_18 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_18 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_18 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_18 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_18 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_18 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_18 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_18 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_18 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_18 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_18 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_18 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_18 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_18 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_18 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_18 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_18 = sboxRom_254;
      default : _zz__zz_stateReg_18 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_7_1)
      8'b00000000 : _zz__zz_stateReg_7 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_7 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_7 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_7 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_7 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_7 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_7 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_7 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_7 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_7 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_7 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_7 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_7 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_7 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_7 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_7 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_7 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_7 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_7 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_7 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_7 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_7 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_7 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_7 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_7 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_7 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_7 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_7 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_7 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_7 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_7 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_7 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_7 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_7 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_7 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_7 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_7 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_7 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_7 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_7 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_7 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_7 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_7 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_7 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_7 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_7 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_7 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_7 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_7 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_7 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_7 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_7 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_7 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_7 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_7 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_7 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_7 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_7 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_7 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_7 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_7 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_7 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_7 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_7 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_7 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_7 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_7 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_7 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_7 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_7 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_7 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_7 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_7 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_7 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_7 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_7 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_7 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_7 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_7 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_7 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_7 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_7 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_7 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_7 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_7 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_7 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_7 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_7 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_7 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_7 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_7 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_7 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_7 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_7 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_7 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_7 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_7 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_7 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_7 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_7 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_7 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_7 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_7 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_7 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_7 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_7 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_7 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_7 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_7 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_7 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_7 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_7 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_7 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_7 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_7 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_7 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_7 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_7 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_7 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_7 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_7 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_7 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_7 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_7 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_7 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_7 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_7 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_7 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_7 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_7 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_7 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_7 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_7 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_7 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_7 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_7 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_7 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_7 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_7 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_7 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_7 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_7 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_7 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_7 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_7 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_7 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_7 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_7 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_7 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_7 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_7 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_7 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_7 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_7 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_7 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_7 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_7 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_7 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_7 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_7 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_7 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_7 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_7 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_7 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_7 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_7 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_7 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_7 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_7 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_7 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_7 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_7 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_7 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_7 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_7 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_7 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_7 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_7 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_7 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_7 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_7 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_7 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_7 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_7 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_7 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_7 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_7 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_7 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_7 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_7 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_7 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_7 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_7 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_7 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_7 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_7 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_7 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_7 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_7 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_7 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_7 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_7 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_7 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_7 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_7 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_7 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_7 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_7 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_7 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_7 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_7 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_7 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_7 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_7 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_7 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_7 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_7 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_7 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_7 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_7 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_7 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_7 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_7 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_7 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_7 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_7 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_7 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_7 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_7 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_7 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_7 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_7 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_7 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_7 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_7 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_7 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_7 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_7 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_7 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_7 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_7 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_7 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_7 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_7 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_7 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_7 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_7 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_7 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_7 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_7 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_7 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_7 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_7 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_7 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_7 = sboxRom_254;
      default : _zz__zz_stateReg_7 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_11_1)
      8'b00000000 : _zz__zz_stateReg_11 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_11 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_11 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_11 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_11 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_11 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_11 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_11 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_11 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_11 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_11 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_11 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_11 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_11 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_11 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_11 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_11 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_11 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_11 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_11 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_11 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_11 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_11 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_11 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_11 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_11 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_11 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_11 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_11 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_11 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_11 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_11 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_11 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_11 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_11 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_11 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_11 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_11 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_11 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_11 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_11 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_11 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_11 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_11 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_11 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_11 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_11 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_11 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_11 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_11 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_11 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_11 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_11 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_11 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_11 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_11 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_11 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_11 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_11 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_11 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_11 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_11 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_11 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_11 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_11 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_11 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_11 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_11 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_11 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_11 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_11 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_11 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_11 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_11 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_11 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_11 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_11 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_11 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_11 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_11 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_11 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_11 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_11 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_11 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_11 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_11 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_11 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_11 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_11 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_11 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_11 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_11 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_11 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_11 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_11 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_11 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_11 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_11 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_11 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_11 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_11 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_11 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_11 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_11 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_11 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_11 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_11 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_11 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_11 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_11 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_11 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_11 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_11 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_11 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_11 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_11 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_11 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_11 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_11 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_11 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_11 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_11 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_11 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_11 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_11 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_11 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_11 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_11 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_11 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_11 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_11 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_11 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_11 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_11 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_11 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_11 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_11 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_11 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_11 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_11 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_11 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_11 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_11 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_11 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_11 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_11 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_11 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_11 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_11 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_11 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_11 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_11 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_11 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_11 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_11 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_11 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_11 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_11 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_11 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_11 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_11 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_11 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_11 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_11 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_11 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_11 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_11 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_11 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_11 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_11 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_11 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_11 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_11 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_11 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_11 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_11 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_11 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_11 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_11 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_11 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_11 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_11 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_11 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_11 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_11 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_11 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_11 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_11 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_11 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_11 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_11 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_11 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_11 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_11 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_11 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_11 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_11 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_11 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_11 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_11 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_11 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_11 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_11 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_11 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_11 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_11 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_11 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_11 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_11 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_11 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_11 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_11 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_11 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_11 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_11 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_11 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_11 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_11 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_11 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_11 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_11 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_11 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_11 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_11 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_11 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_11 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_11 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_11 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_11 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_11 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_11 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_11 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_11 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_11 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_11 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_11 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_11 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_11 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_11 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_11 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_11 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_11 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_11 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_11 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_11 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_11 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_11 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_11 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_11 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_11 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_11 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_11 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_11 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_11 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_11 = sboxRom_254;
      default : _zz__zz_stateReg_11 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_15_1)
      8'b00000000 : _zz__zz_stateReg_15 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_15 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_15 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_15 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_15 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_15 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_15 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_15 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_15 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_15 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_15 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_15 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_15 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_15 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_15 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_15 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_15 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_15 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_15 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_15 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_15 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_15 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_15 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_15 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_15 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_15 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_15 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_15 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_15 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_15 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_15 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_15 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_15 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_15 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_15 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_15 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_15 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_15 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_15 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_15 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_15 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_15 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_15 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_15 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_15 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_15 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_15 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_15 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_15 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_15 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_15 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_15 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_15 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_15 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_15 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_15 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_15 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_15 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_15 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_15 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_15 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_15 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_15 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_15 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_15 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_15 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_15 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_15 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_15 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_15 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_15 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_15 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_15 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_15 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_15 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_15 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_15 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_15 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_15 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_15 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_15 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_15 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_15 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_15 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_15 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_15 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_15 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_15 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_15 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_15 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_15 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_15 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_15 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_15 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_15 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_15 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_15 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_15 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_15 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_15 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_15 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_15 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_15 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_15 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_15 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_15 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_15 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_15 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_15 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_15 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_15 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_15 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_15 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_15 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_15 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_15 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_15 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_15 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_15 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_15 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_15 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_15 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_15 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_15 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_15 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_15 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_15 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_15 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_15 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_15 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_15 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_15 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_15 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_15 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_15 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_15 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_15 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_15 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_15 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_15 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_15 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_15 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_15 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_15 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_15 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_15 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_15 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_15 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_15 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_15 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_15 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_15 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_15 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_15 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_15 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_15 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_15 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_15 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_15 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_15 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_15 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_15 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_15 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_15 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_15 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_15 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_15 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_15 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_15 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_15 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_15 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_15 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_15 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_15 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_15 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_15 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_15 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_15 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_15 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_15 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_15 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_15 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_15 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_15 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_15 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_15 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_15 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_15 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_15 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_15 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_15 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_15 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_15 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_15 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_15 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_15 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_15 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_15 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_15 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_15 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_15 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_15 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_15 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_15 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_15 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_15 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_15 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_15 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_15 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_15 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_15 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_15 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_15 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_15 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_15 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_15 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_15 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_15 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_15 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_15 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_15 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_15 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_15 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_15 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_15 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_15 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_15 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_15 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_15 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_15 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_15 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_15 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_15 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_15 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_15 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_15 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_15 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_15 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_15 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_15 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_15 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_15 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_15 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_15 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_15 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_15 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_15 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_15 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_15 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_15 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_15 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_15 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_15 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_15 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_15 = sboxRom_254;
      default : _zz__zz_stateReg_15 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_19_1)
      8'b00000000 : _zz__zz_stateReg_19 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_19 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_19 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_19 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_19 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_19 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_19 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_19 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_19 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_19 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_19 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_19 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_19 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_19 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_19 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_19 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_19 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_19 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_19 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_19 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_19 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_19 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_19 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_19 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_19 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_19 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_19 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_19 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_19 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_19 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_19 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_19 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_19 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_19 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_19 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_19 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_19 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_19 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_19 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_19 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_19 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_19 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_19 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_19 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_19 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_19 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_19 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_19 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_19 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_19 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_19 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_19 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_19 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_19 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_19 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_19 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_19 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_19 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_19 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_19 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_19 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_19 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_19 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_19 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_19 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_19 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_19 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_19 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_19 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_19 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_19 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_19 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_19 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_19 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_19 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_19 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_19 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_19 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_19 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_19 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_19 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_19 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_19 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_19 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_19 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_19 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_19 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_19 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_19 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_19 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_19 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_19 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_19 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_19 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_19 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_19 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_19 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_19 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_19 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_19 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_19 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_19 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_19 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_19 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_19 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_19 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_19 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_19 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_19 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_19 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_19 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_19 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_19 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_19 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_19 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_19 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_19 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_19 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_19 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_19 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_19 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_19 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_19 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_19 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_19 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_19 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_19 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_19 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_19 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_19 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_19 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_19 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_19 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_19 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_19 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_19 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_19 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_19 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_19 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_19 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_19 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_19 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_19 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_19 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_19 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_19 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_19 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_19 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_19 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_19 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_19 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_19 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_19 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_19 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_19 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_19 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_19 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_19 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_19 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_19 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_19 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_19 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_19 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_19 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_19 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_19 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_19 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_19 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_19 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_19 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_19 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_19 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_19 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_19 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_19 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_19 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_19 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_19 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_19 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_19 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_19 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_19 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_19 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_19 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_19 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_19 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_19 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_19 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_19 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_19 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_19 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_19 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_19 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_19 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_19 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_19 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_19 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_19 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_19 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_19 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_19 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_19 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_19 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_19 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_19 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_19 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_19 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_19 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_19 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_19 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_19 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_19 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_19 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_19 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_19 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_19 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_19 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_19 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_19 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_19 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_19 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_19 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_19 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_19 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_19 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_19 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_19 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_19 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_19 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_19 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_19 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_19 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_19 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_19 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_19 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_19 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_19 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_19 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_19 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_19 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_19 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_19 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_19 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_19 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_19 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_19 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_19 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_19 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_19 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_19 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_19 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_19 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_19 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_19 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_19 = sboxRom_254;
      default : _zz__zz_stateReg_19 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(rconCounter)
      4'b0000 : _zz__zz_roundKeyReg_0 = rcon_0;
      4'b0001 : _zz__zz_roundKeyReg_0 = rcon_1;
      4'b0010 : _zz__zz_roundKeyReg_0 = rcon_2;
      4'b0011 : _zz__zz_roundKeyReg_0 = rcon_3;
      4'b0100 : _zz__zz_roundKeyReg_0 = rcon_4;
      4'b0101 : _zz__zz_roundKeyReg_0 = rcon_5;
      4'b0110 : _zz__zz_roundKeyReg_0 = rcon_6;
      4'b0111 : _zz__zz_roundKeyReg_0 = rcon_7;
      4'b1000 : _zz__zz_roundKeyReg_0 = rcon_8;
      default : _zz__zz_roundKeyReg_0 = rcon_9;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_1)
      8'b00000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_3)
      8'b00000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_5)
      8'b00000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_7)
      8'b00000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_1)
      8'b00000000 : _zz__zz_stateReg_71 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71 = sboxRom_254;
      default : _zz__zz_stateReg_71 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_3)
      8'b00000000 : _zz__zz_stateReg_71_2 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71_2 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71_2 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71_2 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71_2 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71_2 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71_2 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71_2 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71_2 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71_2 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71_2 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71_2 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71_2 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71_2 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71_2 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71_2 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71_2 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71_2 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71_2 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71_2 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71_2 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71_2 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71_2 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71_2 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71_2 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71_2 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71_2 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71_2 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71_2 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71_2 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71_2 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71_2 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71_2 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71_2 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71_2 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71_2 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71_2 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71_2 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71_2 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71_2 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71_2 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71_2 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71_2 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71_2 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71_2 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71_2 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71_2 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71_2 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71_2 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71_2 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71_2 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71_2 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71_2 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71_2 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71_2 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71_2 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71_2 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71_2 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71_2 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71_2 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71_2 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71_2 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71_2 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71_2 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71_2 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71_2 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71_2 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71_2 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71_2 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71_2 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71_2 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71_2 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71_2 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71_2 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71_2 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71_2 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71_2 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71_2 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71_2 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71_2 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71_2 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71_2 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71_2 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71_2 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71_2 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71_2 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71_2 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71_2 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71_2 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71_2 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71_2 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71_2 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71_2 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71_2 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71_2 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71_2 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71_2 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71_2 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71_2 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71_2 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71_2 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71_2 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71_2 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71_2 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71_2 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71_2 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71_2 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71_2 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71_2 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71_2 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71_2 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71_2 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71_2 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71_2 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71_2 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71_2 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71_2 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71_2 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71_2 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71_2 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71_2 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71_2 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71_2 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71_2 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71_2 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71_2 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71_2 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71_2 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71_2 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71_2 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71_2 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71_2 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71_2 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71_2 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71_2 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71_2 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71_2 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71_2 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71_2 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71_2 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71_2 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71_2 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71_2 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71_2 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71_2 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71_2 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71_2 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71_2 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71_2 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71_2 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71_2 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71_2 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71_2 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71_2 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71_2 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71_2 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71_2 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71_2 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71_2 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71_2 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71_2 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71_2 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71_2 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71_2 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71_2 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71_2 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71_2 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71_2 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71_2 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71_2 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71_2 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71_2 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71_2 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71_2 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71_2 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71_2 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71_2 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71_2 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71_2 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71_2 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71_2 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71_2 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71_2 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71_2 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71_2 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71_2 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71_2 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71_2 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71_2 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71_2 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71_2 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71_2 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71_2 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71_2 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71_2 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71_2 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71_2 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71_2 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71_2 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71_2 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71_2 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71_2 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71_2 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71_2 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71_2 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71_2 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71_2 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71_2 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71_2 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71_2 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71_2 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71_2 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71_2 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71_2 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71_2 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71_2 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71_2 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71_2 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71_2 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71_2 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71_2 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71_2 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71_2 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71_2 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71_2 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71_2 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71_2 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71_2 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71_2 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71_2 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71_2 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71_2 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71_2 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71_2 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71_2 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71_2 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71_2 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71_2 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71_2 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71_2 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71_2 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71_2 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71_2 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71_2 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71_2 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71_2 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71_2 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71_2 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71_2 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71_2 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71_2 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71_2 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71_2 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71_2 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71_2 = sboxRom_254;
      default : _zz__zz_stateReg_71_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_5)
      8'b00000000 : _zz__zz_stateReg_71_4 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71_4 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71_4 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71_4 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71_4 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71_4 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71_4 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71_4 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71_4 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71_4 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71_4 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71_4 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71_4 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71_4 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71_4 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71_4 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71_4 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71_4 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71_4 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71_4 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71_4 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71_4 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71_4 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71_4 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71_4 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71_4 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71_4 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71_4 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71_4 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71_4 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71_4 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71_4 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71_4 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71_4 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71_4 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71_4 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71_4 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71_4 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71_4 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71_4 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71_4 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71_4 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71_4 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71_4 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71_4 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71_4 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71_4 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71_4 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71_4 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71_4 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71_4 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71_4 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71_4 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71_4 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71_4 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71_4 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71_4 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71_4 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71_4 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71_4 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71_4 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71_4 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71_4 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71_4 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71_4 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71_4 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71_4 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71_4 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71_4 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71_4 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71_4 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71_4 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71_4 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71_4 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71_4 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71_4 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71_4 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71_4 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71_4 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71_4 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71_4 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71_4 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71_4 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71_4 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71_4 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71_4 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71_4 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71_4 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71_4 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71_4 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71_4 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71_4 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71_4 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71_4 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71_4 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71_4 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71_4 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71_4 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71_4 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71_4 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71_4 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71_4 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71_4 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71_4 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71_4 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71_4 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71_4 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71_4 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71_4 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71_4 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71_4 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71_4 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71_4 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71_4 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71_4 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71_4 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71_4 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71_4 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71_4 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71_4 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71_4 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71_4 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71_4 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71_4 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71_4 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71_4 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71_4 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71_4 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71_4 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71_4 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71_4 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71_4 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71_4 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71_4 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71_4 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71_4 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71_4 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71_4 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71_4 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71_4 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71_4 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71_4 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71_4 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71_4 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71_4 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71_4 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71_4 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71_4 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71_4 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71_4 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71_4 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71_4 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71_4 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71_4 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71_4 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71_4 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71_4 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71_4 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71_4 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71_4 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71_4 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71_4 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71_4 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71_4 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71_4 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71_4 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71_4 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71_4 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71_4 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71_4 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71_4 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71_4 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71_4 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71_4 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71_4 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71_4 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71_4 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71_4 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71_4 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71_4 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71_4 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71_4 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71_4 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71_4 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71_4 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71_4 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71_4 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71_4 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71_4 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71_4 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71_4 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71_4 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71_4 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71_4 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71_4 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71_4 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71_4 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71_4 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71_4 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71_4 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71_4 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71_4 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71_4 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71_4 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71_4 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71_4 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71_4 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71_4 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71_4 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71_4 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71_4 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71_4 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71_4 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71_4 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71_4 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71_4 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71_4 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71_4 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71_4 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71_4 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71_4 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71_4 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71_4 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71_4 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71_4 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71_4 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71_4 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71_4 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71_4 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71_4 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71_4 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71_4 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71_4 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71_4 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71_4 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71_4 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71_4 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71_4 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71_4 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71_4 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71_4 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71_4 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71_4 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71_4 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71_4 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71_4 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71_4 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71_4 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71_4 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71_4 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71_4 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71_4 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71_4 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71_4 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71_4 = sboxRom_254;
      default : _zz__zz_stateReg_71_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_7)
      8'b00000000 : _zz__zz_stateReg_71_6 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71_6 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71_6 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71_6 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71_6 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71_6 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71_6 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71_6 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71_6 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71_6 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71_6 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71_6 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71_6 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71_6 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71_6 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71_6 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71_6 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71_6 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71_6 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71_6 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71_6 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71_6 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71_6 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71_6 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71_6 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71_6 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71_6 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71_6 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71_6 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71_6 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71_6 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71_6 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71_6 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71_6 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71_6 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71_6 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71_6 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71_6 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71_6 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71_6 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71_6 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71_6 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71_6 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71_6 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71_6 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71_6 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71_6 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71_6 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71_6 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71_6 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71_6 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71_6 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71_6 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71_6 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71_6 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71_6 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71_6 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71_6 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71_6 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71_6 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71_6 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71_6 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71_6 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71_6 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71_6 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71_6 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71_6 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71_6 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71_6 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71_6 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71_6 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71_6 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71_6 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71_6 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71_6 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71_6 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71_6 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71_6 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71_6 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71_6 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71_6 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71_6 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71_6 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71_6 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71_6 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71_6 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71_6 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71_6 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71_6 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71_6 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71_6 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71_6 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71_6 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71_6 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71_6 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71_6 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71_6 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71_6 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71_6 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71_6 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71_6 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71_6 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71_6 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71_6 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71_6 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71_6 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71_6 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71_6 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71_6 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71_6 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71_6 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71_6 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71_6 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71_6 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71_6 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71_6 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71_6 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71_6 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71_6 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71_6 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71_6 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71_6 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71_6 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71_6 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71_6 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71_6 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71_6 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71_6 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71_6 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71_6 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71_6 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71_6 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71_6 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71_6 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71_6 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71_6 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71_6 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71_6 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71_6 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71_6 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71_6 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71_6 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71_6 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71_6 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71_6 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71_6 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71_6 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71_6 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71_6 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71_6 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71_6 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71_6 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71_6 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71_6 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71_6 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71_6 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71_6 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71_6 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71_6 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71_6 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71_6 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71_6 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71_6 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71_6 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71_6 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71_6 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71_6 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71_6 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71_6 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71_6 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71_6 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71_6 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71_6 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71_6 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71_6 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71_6 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71_6 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71_6 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71_6 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71_6 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71_6 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71_6 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71_6 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71_6 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71_6 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71_6 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71_6 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71_6 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71_6 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71_6 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71_6 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71_6 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71_6 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71_6 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71_6 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71_6 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71_6 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71_6 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71_6 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71_6 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71_6 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71_6 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71_6 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71_6 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71_6 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71_6 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71_6 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71_6 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71_6 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71_6 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71_6 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71_6 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71_6 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71_6 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71_6 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71_6 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71_6 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71_6 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71_6 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71_6 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71_6 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71_6 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71_6 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71_6 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71_6 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71_6 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71_6 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71_6 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71_6 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71_6 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71_6 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71_6 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71_6 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71_6 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71_6 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71_6 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71_6 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71_6 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71_6 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71_6 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71_6 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71_6 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71_6 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71_6 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71_6 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71_6 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71_6 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71_6 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71_6 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71_6 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71_6 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71_6 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71_6 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71_6 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71_6 = sboxRom_254;
      default : _zz__zz_stateReg_71_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(precomputeCounter)
      4'b0000 : _zz__zz_stateReg_71_8 = rcon_0;
      4'b0001 : _zz__zz_stateReg_71_8 = rcon_1;
      4'b0010 : _zz__zz_stateReg_71_8 = rcon_2;
      4'b0011 : _zz__zz_stateReg_71_8 = rcon_3;
      4'b0100 : _zz__zz_stateReg_71_8 = rcon_4;
      4'b0101 : _zz__zz_stateReg_71_8 = rcon_5;
      4'b0110 : _zz__zz_stateReg_71_8 = rcon_6;
      4'b0111 : _zz__zz_stateReg_71_8 = rcon_7;
      4'b1000 : _zz__zz_stateReg_71_8 = rcon_8;
      default : _zz__zz_stateReg_71_8 = rcon_9;
    endcase
  end

  always @(*) begin
    case(invShifted_0)
      8'b00000000 : _zz_invSub_0 = invSboxRom_0;
      8'b00000001 : _zz_invSub_0 = invSboxRom_1;
      8'b00000010 : _zz_invSub_0 = invSboxRom_2;
      8'b00000011 : _zz_invSub_0 = invSboxRom_3;
      8'b00000100 : _zz_invSub_0 = invSboxRom_4;
      8'b00000101 : _zz_invSub_0 = invSboxRom_5;
      8'b00000110 : _zz_invSub_0 = invSboxRom_6;
      8'b00000111 : _zz_invSub_0 = invSboxRom_7;
      8'b00001000 : _zz_invSub_0 = invSboxRom_8;
      8'b00001001 : _zz_invSub_0 = invSboxRom_9;
      8'b00001010 : _zz_invSub_0 = invSboxRom_10;
      8'b00001011 : _zz_invSub_0 = invSboxRom_11;
      8'b00001100 : _zz_invSub_0 = invSboxRom_12;
      8'b00001101 : _zz_invSub_0 = invSboxRom_13;
      8'b00001110 : _zz_invSub_0 = invSboxRom_14;
      8'b00001111 : _zz_invSub_0 = invSboxRom_15;
      8'b00010000 : _zz_invSub_0 = invSboxRom_16;
      8'b00010001 : _zz_invSub_0 = invSboxRom_17;
      8'b00010010 : _zz_invSub_0 = invSboxRom_18;
      8'b00010011 : _zz_invSub_0 = invSboxRom_19;
      8'b00010100 : _zz_invSub_0 = invSboxRom_20;
      8'b00010101 : _zz_invSub_0 = invSboxRom_21;
      8'b00010110 : _zz_invSub_0 = invSboxRom_22;
      8'b00010111 : _zz_invSub_0 = invSboxRom_23;
      8'b00011000 : _zz_invSub_0 = invSboxRom_24;
      8'b00011001 : _zz_invSub_0 = invSboxRom_25;
      8'b00011010 : _zz_invSub_0 = invSboxRom_26;
      8'b00011011 : _zz_invSub_0 = invSboxRom_27;
      8'b00011100 : _zz_invSub_0 = invSboxRom_28;
      8'b00011101 : _zz_invSub_0 = invSboxRom_29;
      8'b00011110 : _zz_invSub_0 = invSboxRom_30;
      8'b00011111 : _zz_invSub_0 = invSboxRom_31;
      8'b00100000 : _zz_invSub_0 = invSboxRom_32;
      8'b00100001 : _zz_invSub_0 = invSboxRom_33;
      8'b00100010 : _zz_invSub_0 = invSboxRom_34;
      8'b00100011 : _zz_invSub_0 = invSboxRom_35;
      8'b00100100 : _zz_invSub_0 = invSboxRom_36;
      8'b00100101 : _zz_invSub_0 = invSboxRom_37;
      8'b00100110 : _zz_invSub_0 = invSboxRom_38;
      8'b00100111 : _zz_invSub_0 = invSboxRom_39;
      8'b00101000 : _zz_invSub_0 = invSboxRom_40;
      8'b00101001 : _zz_invSub_0 = invSboxRom_41;
      8'b00101010 : _zz_invSub_0 = invSboxRom_42;
      8'b00101011 : _zz_invSub_0 = invSboxRom_43;
      8'b00101100 : _zz_invSub_0 = invSboxRom_44;
      8'b00101101 : _zz_invSub_0 = invSboxRom_45;
      8'b00101110 : _zz_invSub_0 = invSboxRom_46;
      8'b00101111 : _zz_invSub_0 = invSboxRom_47;
      8'b00110000 : _zz_invSub_0 = invSboxRom_48;
      8'b00110001 : _zz_invSub_0 = invSboxRom_49;
      8'b00110010 : _zz_invSub_0 = invSboxRom_50;
      8'b00110011 : _zz_invSub_0 = invSboxRom_51;
      8'b00110100 : _zz_invSub_0 = invSboxRom_52;
      8'b00110101 : _zz_invSub_0 = invSboxRom_53;
      8'b00110110 : _zz_invSub_0 = invSboxRom_54;
      8'b00110111 : _zz_invSub_0 = invSboxRom_55;
      8'b00111000 : _zz_invSub_0 = invSboxRom_56;
      8'b00111001 : _zz_invSub_0 = invSboxRom_57;
      8'b00111010 : _zz_invSub_0 = invSboxRom_58;
      8'b00111011 : _zz_invSub_0 = invSboxRom_59;
      8'b00111100 : _zz_invSub_0 = invSboxRom_60;
      8'b00111101 : _zz_invSub_0 = invSboxRom_61;
      8'b00111110 : _zz_invSub_0 = invSboxRom_62;
      8'b00111111 : _zz_invSub_0 = invSboxRom_63;
      8'b01000000 : _zz_invSub_0 = invSboxRom_64;
      8'b01000001 : _zz_invSub_0 = invSboxRom_65;
      8'b01000010 : _zz_invSub_0 = invSboxRom_66;
      8'b01000011 : _zz_invSub_0 = invSboxRom_67;
      8'b01000100 : _zz_invSub_0 = invSboxRom_68;
      8'b01000101 : _zz_invSub_0 = invSboxRom_69;
      8'b01000110 : _zz_invSub_0 = invSboxRom_70;
      8'b01000111 : _zz_invSub_0 = invSboxRom_71;
      8'b01001000 : _zz_invSub_0 = invSboxRom_72;
      8'b01001001 : _zz_invSub_0 = invSboxRom_73;
      8'b01001010 : _zz_invSub_0 = invSboxRom_74;
      8'b01001011 : _zz_invSub_0 = invSboxRom_75;
      8'b01001100 : _zz_invSub_0 = invSboxRom_76;
      8'b01001101 : _zz_invSub_0 = invSboxRom_77;
      8'b01001110 : _zz_invSub_0 = invSboxRom_78;
      8'b01001111 : _zz_invSub_0 = invSboxRom_79;
      8'b01010000 : _zz_invSub_0 = invSboxRom_80;
      8'b01010001 : _zz_invSub_0 = invSboxRom_81;
      8'b01010010 : _zz_invSub_0 = invSboxRom_82;
      8'b01010011 : _zz_invSub_0 = invSboxRom_83;
      8'b01010100 : _zz_invSub_0 = invSboxRom_84;
      8'b01010101 : _zz_invSub_0 = invSboxRom_85;
      8'b01010110 : _zz_invSub_0 = invSboxRom_86;
      8'b01010111 : _zz_invSub_0 = invSboxRom_87;
      8'b01011000 : _zz_invSub_0 = invSboxRom_88;
      8'b01011001 : _zz_invSub_0 = invSboxRom_89;
      8'b01011010 : _zz_invSub_0 = invSboxRom_90;
      8'b01011011 : _zz_invSub_0 = invSboxRom_91;
      8'b01011100 : _zz_invSub_0 = invSboxRom_92;
      8'b01011101 : _zz_invSub_0 = invSboxRom_93;
      8'b01011110 : _zz_invSub_0 = invSboxRom_94;
      8'b01011111 : _zz_invSub_0 = invSboxRom_95;
      8'b01100000 : _zz_invSub_0 = invSboxRom_96;
      8'b01100001 : _zz_invSub_0 = invSboxRom_97;
      8'b01100010 : _zz_invSub_0 = invSboxRom_98;
      8'b01100011 : _zz_invSub_0 = invSboxRom_99;
      8'b01100100 : _zz_invSub_0 = invSboxRom_100;
      8'b01100101 : _zz_invSub_0 = invSboxRom_101;
      8'b01100110 : _zz_invSub_0 = invSboxRom_102;
      8'b01100111 : _zz_invSub_0 = invSboxRom_103;
      8'b01101000 : _zz_invSub_0 = invSboxRom_104;
      8'b01101001 : _zz_invSub_0 = invSboxRom_105;
      8'b01101010 : _zz_invSub_0 = invSboxRom_106;
      8'b01101011 : _zz_invSub_0 = invSboxRom_107;
      8'b01101100 : _zz_invSub_0 = invSboxRom_108;
      8'b01101101 : _zz_invSub_0 = invSboxRom_109;
      8'b01101110 : _zz_invSub_0 = invSboxRom_110;
      8'b01101111 : _zz_invSub_0 = invSboxRom_111;
      8'b01110000 : _zz_invSub_0 = invSboxRom_112;
      8'b01110001 : _zz_invSub_0 = invSboxRom_113;
      8'b01110010 : _zz_invSub_0 = invSboxRom_114;
      8'b01110011 : _zz_invSub_0 = invSboxRom_115;
      8'b01110100 : _zz_invSub_0 = invSboxRom_116;
      8'b01110101 : _zz_invSub_0 = invSboxRom_117;
      8'b01110110 : _zz_invSub_0 = invSboxRom_118;
      8'b01110111 : _zz_invSub_0 = invSboxRom_119;
      8'b01111000 : _zz_invSub_0 = invSboxRom_120;
      8'b01111001 : _zz_invSub_0 = invSboxRom_121;
      8'b01111010 : _zz_invSub_0 = invSboxRom_122;
      8'b01111011 : _zz_invSub_0 = invSboxRom_123;
      8'b01111100 : _zz_invSub_0 = invSboxRom_124;
      8'b01111101 : _zz_invSub_0 = invSboxRom_125;
      8'b01111110 : _zz_invSub_0 = invSboxRom_126;
      8'b01111111 : _zz_invSub_0 = invSboxRom_127;
      8'b10000000 : _zz_invSub_0 = invSboxRom_128;
      8'b10000001 : _zz_invSub_0 = invSboxRom_129;
      8'b10000010 : _zz_invSub_0 = invSboxRom_130;
      8'b10000011 : _zz_invSub_0 = invSboxRom_131;
      8'b10000100 : _zz_invSub_0 = invSboxRom_132;
      8'b10000101 : _zz_invSub_0 = invSboxRom_133;
      8'b10000110 : _zz_invSub_0 = invSboxRom_134;
      8'b10000111 : _zz_invSub_0 = invSboxRom_135;
      8'b10001000 : _zz_invSub_0 = invSboxRom_136;
      8'b10001001 : _zz_invSub_0 = invSboxRom_137;
      8'b10001010 : _zz_invSub_0 = invSboxRom_138;
      8'b10001011 : _zz_invSub_0 = invSboxRom_139;
      8'b10001100 : _zz_invSub_0 = invSboxRom_140;
      8'b10001101 : _zz_invSub_0 = invSboxRom_141;
      8'b10001110 : _zz_invSub_0 = invSboxRom_142;
      8'b10001111 : _zz_invSub_0 = invSboxRom_143;
      8'b10010000 : _zz_invSub_0 = invSboxRom_144;
      8'b10010001 : _zz_invSub_0 = invSboxRom_145;
      8'b10010010 : _zz_invSub_0 = invSboxRom_146;
      8'b10010011 : _zz_invSub_0 = invSboxRom_147;
      8'b10010100 : _zz_invSub_0 = invSboxRom_148;
      8'b10010101 : _zz_invSub_0 = invSboxRom_149;
      8'b10010110 : _zz_invSub_0 = invSboxRom_150;
      8'b10010111 : _zz_invSub_0 = invSboxRom_151;
      8'b10011000 : _zz_invSub_0 = invSboxRom_152;
      8'b10011001 : _zz_invSub_0 = invSboxRom_153;
      8'b10011010 : _zz_invSub_0 = invSboxRom_154;
      8'b10011011 : _zz_invSub_0 = invSboxRom_155;
      8'b10011100 : _zz_invSub_0 = invSboxRom_156;
      8'b10011101 : _zz_invSub_0 = invSboxRom_157;
      8'b10011110 : _zz_invSub_0 = invSboxRom_158;
      8'b10011111 : _zz_invSub_0 = invSboxRom_159;
      8'b10100000 : _zz_invSub_0 = invSboxRom_160;
      8'b10100001 : _zz_invSub_0 = invSboxRom_161;
      8'b10100010 : _zz_invSub_0 = invSboxRom_162;
      8'b10100011 : _zz_invSub_0 = invSboxRom_163;
      8'b10100100 : _zz_invSub_0 = invSboxRom_164;
      8'b10100101 : _zz_invSub_0 = invSboxRom_165;
      8'b10100110 : _zz_invSub_0 = invSboxRom_166;
      8'b10100111 : _zz_invSub_0 = invSboxRom_167;
      8'b10101000 : _zz_invSub_0 = invSboxRom_168;
      8'b10101001 : _zz_invSub_0 = invSboxRom_169;
      8'b10101010 : _zz_invSub_0 = invSboxRom_170;
      8'b10101011 : _zz_invSub_0 = invSboxRom_171;
      8'b10101100 : _zz_invSub_0 = invSboxRom_172;
      8'b10101101 : _zz_invSub_0 = invSboxRom_173;
      8'b10101110 : _zz_invSub_0 = invSboxRom_174;
      8'b10101111 : _zz_invSub_0 = invSboxRom_175;
      8'b10110000 : _zz_invSub_0 = invSboxRom_176;
      8'b10110001 : _zz_invSub_0 = invSboxRom_177;
      8'b10110010 : _zz_invSub_0 = invSboxRom_178;
      8'b10110011 : _zz_invSub_0 = invSboxRom_179;
      8'b10110100 : _zz_invSub_0 = invSboxRom_180;
      8'b10110101 : _zz_invSub_0 = invSboxRom_181;
      8'b10110110 : _zz_invSub_0 = invSboxRom_182;
      8'b10110111 : _zz_invSub_0 = invSboxRom_183;
      8'b10111000 : _zz_invSub_0 = invSboxRom_184;
      8'b10111001 : _zz_invSub_0 = invSboxRom_185;
      8'b10111010 : _zz_invSub_0 = invSboxRom_186;
      8'b10111011 : _zz_invSub_0 = invSboxRom_187;
      8'b10111100 : _zz_invSub_0 = invSboxRom_188;
      8'b10111101 : _zz_invSub_0 = invSboxRom_189;
      8'b10111110 : _zz_invSub_0 = invSboxRom_190;
      8'b10111111 : _zz_invSub_0 = invSboxRom_191;
      8'b11000000 : _zz_invSub_0 = invSboxRom_192;
      8'b11000001 : _zz_invSub_0 = invSboxRom_193;
      8'b11000010 : _zz_invSub_0 = invSboxRom_194;
      8'b11000011 : _zz_invSub_0 = invSboxRom_195;
      8'b11000100 : _zz_invSub_0 = invSboxRom_196;
      8'b11000101 : _zz_invSub_0 = invSboxRom_197;
      8'b11000110 : _zz_invSub_0 = invSboxRom_198;
      8'b11000111 : _zz_invSub_0 = invSboxRom_199;
      8'b11001000 : _zz_invSub_0 = invSboxRom_200;
      8'b11001001 : _zz_invSub_0 = invSboxRom_201;
      8'b11001010 : _zz_invSub_0 = invSboxRom_202;
      8'b11001011 : _zz_invSub_0 = invSboxRom_203;
      8'b11001100 : _zz_invSub_0 = invSboxRom_204;
      8'b11001101 : _zz_invSub_0 = invSboxRom_205;
      8'b11001110 : _zz_invSub_0 = invSboxRom_206;
      8'b11001111 : _zz_invSub_0 = invSboxRom_207;
      8'b11010000 : _zz_invSub_0 = invSboxRom_208;
      8'b11010001 : _zz_invSub_0 = invSboxRom_209;
      8'b11010010 : _zz_invSub_0 = invSboxRom_210;
      8'b11010011 : _zz_invSub_0 = invSboxRom_211;
      8'b11010100 : _zz_invSub_0 = invSboxRom_212;
      8'b11010101 : _zz_invSub_0 = invSboxRom_213;
      8'b11010110 : _zz_invSub_0 = invSboxRom_214;
      8'b11010111 : _zz_invSub_0 = invSboxRom_215;
      8'b11011000 : _zz_invSub_0 = invSboxRom_216;
      8'b11011001 : _zz_invSub_0 = invSboxRom_217;
      8'b11011010 : _zz_invSub_0 = invSboxRom_218;
      8'b11011011 : _zz_invSub_0 = invSboxRom_219;
      8'b11011100 : _zz_invSub_0 = invSboxRom_220;
      8'b11011101 : _zz_invSub_0 = invSboxRom_221;
      8'b11011110 : _zz_invSub_0 = invSboxRom_222;
      8'b11011111 : _zz_invSub_0 = invSboxRom_223;
      8'b11100000 : _zz_invSub_0 = invSboxRom_224;
      8'b11100001 : _zz_invSub_0 = invSboxRom_225;
      8'b11100010 : _zz_invSub_0 = invSboxRom_226;
      8'b11100011 : _zz_invSub_0 = invSboxRom_227;
      8'b11100100 : _zz_invSub_0 = invSboxRom_228;
      8'b11100101 : _zz_invSub_0 = invSboxRom_229;
      8'b11100110 : _zz_invSub_0 = invSboxRom_230;
      8'b11100111 : _zz_invSub_0 = invSboxRom_231;
      8'b11101000 : _zz_invSub_0 = invSboxRom_232;
      8'b11101001 : _zz_invSub_0 = invSboxRom_233;
      8'b11101010 : _zz_invSub_0 = invSboxRom_234;
      8'b11101011 : _zz_invSub_0 = invSboxRom_235;
      8'b11101100 : _zz_invSub_0 = invSboxRom_236;
      8'b11101101 : _zz_invSub_0 = invSboxRom_237;
      8'b11101110 : _zz_invSub_0 = invSboxRom_238;
      8'b11101111 : _zz_invSub_0 = invSboxRom_239;
      8'b11110000 : _zz_invSub_0 = invSboxRom_240;
      8'b11110001 : _zz_invSub_0 = invSboxRom_241;
      8'b11110010 : _zz_invSub_0 = invSboxRom_242;
      8'b11110011 : _zz_invSub_0 = invSboxRom_243;
      8'b11110100 : _zz_invSub_0 = invSboxRom_244;
      8'b11110101 : _zz_invSub_0 = invSboxRom_245;
      8'b11110110 : _zz_invSub_0 = invSboxRom_246;
      8'b11110111 : _zz_invSub_0 = invSboxRom_247;
      8'b11111000 : _zz_invSub_0 = invSboxRom_248;
      8'b11111001 : _zz_invSub_0 = invSboxRom_249;
      8'b11111010 : _zz_invSub_0 = invSboxRom_250;
      8'b11111011 : _zz_invSub_0 = invSboxRom_251;
      8'b11111100 : _zz_invSub_0 = invSboxRom_252;
      8'b11111101 : _zz_invSub_0 = invSboxRom_253;
      8'b11111110 : _zz_invSub_0 = invSboxRom_254;
      default : _zz_invSub_0 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_1)
      8'b00000000 : _zz_invSub_1 = invSboxRom_0;
      8'b00000001 : _zz_invSub_1 = invSboxRom_1;
      8'b00000010 : _zz_invSub_1 = invSboxRom_2;
      8'b00000011 : _zz_invSub_1 = invSboxRom_3;
      8'b00000100 : _zz_invSub_1 = invSboxRom_4;
      8'b00000101 : _zz_invSub_1 = invSboxRom_5;
      8'b00000110 : _zz_invSub_1 = invSboxRom_6;
      8'b00000111 : _zz_invSub_1 = invSboxRom_7;
      8'b00001000 : _zz_invSub_1 = invSboxRom_8;
      8'b00001001 : _zz_invSub_1 = invSboxRom_9;
      8'b00001010 : _zz_invSub_1 = invSboxRom_10;
      8'b00001011 : _zz_invSub_1 = invSboxRom_11;
      8'b00001100 : _zz_invSub_1 = invSboxRom_12;
      8'b00001101 : _zz_invSub_1 = invSboxRom_13;
      8'b00001110 : _zz_invSub_1 = invSboxRom_14;
      8'b00001111 : _zz_invSub_1 = invSboxRom_15;
      8'b00010000 : _zz_invSub_1 = invSboxRom_16;
      8'b00010001 : _zz_invSub_1 = invSboxRom_17;
      8'b00010010 : _zz_invSub_1 = invSboxRom_18;
      8'b00010011 : _zz_invSub_1 = invSboxRom_19;
      8'b00010100 : _zz_invSub_1 = invSboxRom_20;
      8'b00010101 : _zz_invSub_1 = invSboxRom_21;
      8'b00010110 : _zz_invSub_1 = invSboxRom_22;
      8'b00010111 : _zz_invSub_1 = invSboxRom_23;
      8'b00011000 : _zz_invSub_1 = invSboxRom_24;
      8'b00011001 : _zz_invSub_1 = invSboxRom_25;
      8'b00011010 : _zz_invSub_1 = invSboxRom_26;
      8'b00011011 : _zz_invSub_1 = invSboxRom_27;
      8'b00011100 : _zz_invSub_1 = invSboxRom_28;
      8'b00011101 : _zz_invSub_1 = invSboxRom_29;
      8'b00011110 : _zz_invSub_1 = invSboxRom_30;
      8'b00011111 : _zz_invSub_1 = invSboxRom_31;
      8'b00100000 : _zz_invSub_1 = invSboxRom_32;
      8'b00100001 : _zz_invSub_1 = invSboxRom_33;
      8'b00100010 : _zz_invSub_1 = invSboxRom_34;
      8'b00100011 : _zz_invSub_1 = invSboxRom_35;
      8'b00100100 : _zz_invSub_1 = invSboxRom_36;
      8'b00100101 : _zz_invSub_1 = invSboxRom_37;
      8'b00100110 : _zz_invSub_1 = invSboxRom_38;
      8'b00100111 : _zz_invSub_1 = invSboxRom_39;
      8'b00101000 : _zz_invSub_1 = invSboxRom_40;
      8'b00101001 : _zz_invSub_1 = invSboxRom_41;
      8'b00101010 : _zz_invSub_1 = invSboxRom_42;
      8'b00101011 : _zz_invSub_1 = invSboxRom_43;
      8'b00101100 : _zz_invSub_1 = invSboxRom_44;
      8'b00101101 : _zz_invSub_1 = invSboxRom_45;
      8'b00101110 : _zz_invSub_1 = invSboxRom_46;
      8'b00101111 : _zz_invSub_1 = invSboxRom_47;
      8'b00110000 : _zz_invSub_1 = invSboxRom_48;
      8'b00110001 : _zz_invSub_1 = invSboxRom_49;
      8'b00110010 : _zz_invSub_1 = invSboxRom_50;
      8'b00110011 : _zz_invSub_1 = invSboxRom_51;
      8'b00110100 : _zz_invSub_1 = invSboxRom_52;
      8'b00110101 : _zz_invSub_1 = invSboxRom_53;
      8'b00110110 : _zz_invSub_1 = invSboxRom_54;
      8'b00110111 : _zz_invSub_1 = invSboxRom_55;
      8'b00111000 : _zz_invSub_1 = invSboxRom_56;
      8'b00111001 : _zz_invSub_1 = invSboxRom_57;
      8'b00111010 : _zz_invSub_1 = invSboxRom_58;
      8'b00111011 : _zz_invSub_1 = invSboxRom_59;
      8'b00111100 : _zz_invSub_1 = invSboxRom_60;
      8'b00111101 : _zz_invSub_1 = invSboxRom_61;
      8'b00111110 : _zz_invSub_1 = invSboxRom_62;
      8'b00111111 : _zz_invSub_1 = invSboxRom_63;
      8'b01000000 : _zz_invSub_1 = invSboxRom_64;
      8'b01000001 : _zz_invSub_1 = invSboxRom_65;
      8'b01000010 : _zz_invSub_1 = invSboxRom_66;
      8'b01000011 : _zz_invSub_1 = invSboxRom_67;
      8'b01000100 : _zz_invSub_1 = invSboxRom_68;
      8'b01000101 : _zz_invSub_1 = invSboxRom_69;
      8'b01000110 : _zz_invSub_1 = invSboxRom_70;
      8'b01000111 : _zz_invSub_1 = invSboxRom_71;
      8'b01001000 : _zz_invSub_1 = invSboxRom_72;
      8'b01001001 : _zz_invSub_1 = invSboxRom_73;
      8'b01001010 : _zz_invSub_1 = invSboxRom_74;
      8'b01001011 : _zz_invSub_1 = invSboxRom_75;
      8'b01001100 : _zz_invSub_1 = invSboxRom_76;
      8'b01001101 : _zz_invSub_1 = invSboxRom_77;
      8'b01001110 : _zz_invSub_1 = invSboxRom_78;
      8'b01001111 : _zz_invSub_1 = invSboxRom_79;
      8'b01010000 : _zz_invSub_1 = invSboxRom_80;
      8'b01010001 : _zz_invSub_1 = invSboxRom_81;
      8'b01010010 : _zz_invSub_1 = invSboxRom_82;
      8'b01010011 : _zz_invSub_1 = invSboxRom_83;
      8'b01010100 : _zz_invSub_1 = invSboxRom_84;
      8'b01010101 : _zz_invSub_1 = invSboxRom_85;
      8'b01010110 : _zz_invSub_1 = invSboxRom_86;
      8'b01010111 : _zz_invSub_1 = invSboxRom_87;
      8'b01011000 : _zz_invSub_1 = invSboxRom_88;
      8'b01011001 : _zz_invSub_1 = invSboxRom_89;
      8'b01011010 : _zz_invSub_1 = invSboxRom_90;
      8'b01011011 : _zz_invSub_1 = invSboxRom_91;
      8'b01011100 : _zz_invSub_1 = invSboxRom_92;
      8'b01011101 : _zz_invSub_1 = invSboxRom_93;
      8'b01011110 : _zz_invSub_1 = invSboxRom_94;
      8'b01011111 : _zz_invSub_1 = invSboxRom_95;
      8'b01100000 : _zz_invSub_1 = invSboxRom_96;
      8'b01100001 : _zz_invSub_1 = invSboxRom_97;
      8'b01100010 : _zz_invSub_1 = invSboxRom_98;
      8'b01100011 : _zz_invSub_1 = invSboxRom_99;
      8'b01100100 : _zz_invSub_1 = invSboxRom_100;
      8'b01100101 : _zz_invSub_1 = invSboxRom_101;
      8'b01100110 : _zz_invSub_1 = invSboxRom_102;
      8'b01100111 : _zz_invSub_1 = invSboxRom_103;
      8'b01101000 : _zz_invSub_1 = invSboxRom_104;
      8'b01101001 : _zz_invSub_1 = invSboxRom_105;
      8'b01101010 : _zz_invSub_1 = invSboxRom_106;
      8'b01101011 : _zz_invSub_1 = invSboxRom_107;
      8'b01101100 : _zz_invSub_1 = invSboxRom_108;
      8'b01101101 : _zz_invSub_1 = invSboxRom_109;
      8'b01101110 : _zz_invSub_1 = invSboxRom_110;
      8'b01101111 : _zz_invSub_1 = invSboxRom_111;
      8'b01110000 : _zz_invSub_1 = invSboxRom_112;
      8'b01110001 : _zz_invSub_1 = invSboxRom_113;
      8'b01110010 : _zz_invSub_1 = invSboxRom_114;
      8'b01110011 : _zz_invSub_1 = invSboxRom_115;
      8'b01110100 : _zz_invSub_1 = invSboxRom_116;
      8'b01110101 : _zz_invSub_1 = invSboxRom_117;
      8'b01110110 : _zz_invSub_1 = invSboxRom_118;
      8'b01110111 : _zz_invSub_1 = invSboxRom_119;
      8'b01111000 : _zz_invSub_1 = invSboxRom_120;
      8'b01111001 : _zz_invSub_1 = invSboxRom_121;
      8'b01111010 : _zz_invSub_1 = invSboxRom_122;
      8'b01111011 : _zz_invSub_1 = invSboxRom_123;
      8'b01111100 : _zz_invSub_1 = invSboxRom_124;
      8'b01111101 : _zz_invSub_1 = invSboxRom_125;
      8'b01111110 : _zz_invSub_1 = invSboxRom_126;
      8'b01111111 : _zz_invSub_1 = invSboxRom_127;
      8'b10000000 : _zz_invSub_1 = invSboxRom_128;
      8'b10000001 : _zz_invSub_1 = invSboxRom_129;
      8'b10000010 : _zz_invSub_1 = invSboxRom_130;
      8'b10000011 : _zz_invSub_1 = invSboxRom_131;
      8'b10000100 : _zz_invSub_1 = invSboxRom_132;
      8'b10000101 : _zz_invSub_1 = invSboxRom_133;
      8'b10000110 : _zz_invSub_1 = invSboxRom_134;
      8'b10000111 : _zz_invSub_1 = invSboxRom_135;
      8'b10001000 : _zz_invSub_1 = invSboxRom_136;
      8'b10001001 : _zz_invSub_1 = invSboxRom_137;
      8'b10001010 : _zz_invSub_1 = invSboxRom_138;
      8'b10001011 : _zz_invSub_1 = invSboxRom_139;
      8'b10001100 : _zz_invSub_1 = invSboxRom_140;
      8'b10001101 : _zz_invSub_1 = invSboxRom_141;
      8'b10001110 : _zz_invSub_1 = invSboxRom_142;
      8'b10001111 : _zz_invSub_1 = invSboxRom_143;
      8'b10010000 : _zz_invSub_1 = invSboxRom_144;
      8'b10010001 : _zz_invSub_1 = invSboxRom_145;
      8'b10010010 : _zz_invSub_1 = invSboxRom_146;
      8'b10010011 : _zz_invSub_1 = invSboxRom_147;
      8'b10010100 : _zz_invSub_1 = invSboxRom_148;
      8'b10010101 : _zz_invSub_1 = invSboxRom_149;
      8'b10010110 : _zz_invSub_1 = invSboxRom_150;
      8'b10010111 : _zz_invSub_1 = invSboxRom_151;
      8'b10011000 : _zz_invSub_1 = invSboxRom_152;
      8'b10011001 : _zz_invSub_1 = invSboxRom_153;
      8'b10011010 : _zz_invSub_1 = invSboxRom_154;
      8'b10011011 : _zz_invSub_1 = invSboxRom_155;
      8'b10011100 : _zz_invSub_1 = invSboxRom_156;
      8'b10011101 : _zz_invSub_1 = invSboxRom_157;
      8'b10011110 : _zz_invSub_1 = invSboxRom_158;
      8'b10011111 : _zz_invSub_1 = invSboxRom_159;
      8'b10100000 : _zz_invSub_1 = invSboxRom_160;
      8'b10100001 : _zz_invSub_1 = invSboxRom_161;
      8'b10100010 : _zz_invSub_1 = invSboxRom_162;
      8'b10100011 : _zz_invSub_1 = invSboxRom_163;
      8'b10100100 : _zz_invSub_1 = invSboxRom_164;
      8'b10100101 : _zz_invSub_1 = invSboxRom_165;
      8'b10100110 : _zz_invSub_1 = invSboxRom_166;
      8'b10100111 : _zz_invSub_1 = invSboxRom_167;
      8'b10101000 : _zz_invSub_1 = invSboxRom_168;
      8'b10101001 : _zz_invSub_1 = invSboxRom_169;
      8'b10101010 : _zz_invSub_1 = invSboxRom_170;
      8'b10101011 : _zz_invSub_1 = invSboxRom_171;
      8'b10101100 : _zz_invSub_1 = invSboxRom_172;
      8'b10101101 : _zz_invSub_1 = invSboxRom_173;
      8'b10101110 : _zz_invSub_1 = invSboxRom_174;
      8'b10101111 : _zz_invSub_1 = invSboxRom_175;
      8'b10110000 : _zz_invSub_1 = invSboxRom_176;
      8'b10110001 : _zz_invSub_1 = invSboxRom_177;
      8'b10110010 : _zz_invSub_1 = invSboxRom_178;
      8'b10110011 : _zz_invSub_1 = invSboxRom_179;
      8'b10110100 : _zz_invSub_1 = invSboxRom_180;
      8'b10110101 : _zz_invSub_1 = invSboxRom_181;
      8'b10110110 : _zz_invSub_1 = invSboxRom_182;
      8'b10110111 : _zz_invSub_1 = invSboxRom_183;
      8'b10111000 : _zz_invSub_1 = invSboxRom_184;
      8'b10111001 : _zz_invSub_1 = invSboxRom_185;
      8'b10111010 : _zz_invSub_1 = invSboxRom_186;
      8'b10111011 : _zz_invSub_1 = invSboxRom_187;
      8'b10111100 : _zz_invSub_1 = invSboxRom_188;
      8'b10111101 : _zz_invSub_1 = invSboxRom_189;
      8'b10111110 : _zz_invSub_1 = invSboxRom_190;
      8'b10111111 : _zz_invSub_1 = invSboxRom_191;
      8'b11000000 : _zz_invSub_1 = invSboxRom_192;
      8'b11000001 : _zz_invSub_1 = invSboxRom_193;
      8'b11000010 : _zz_invSub_1 = invSboxRom_194;
      8'b11000011 : _zz_invSub_1 = invSboxRom_195;
      8'b11000100 : _zz_invSub_1 = invSboxRom_196;
      8'b11000101 : _zz_invSub_1 = invSboxRom_197;
      8'b11000110 : _zz_invSub_1 = invSboxRom_198;
      8'b11000111 : _zz_invSub_1 = invSboxRom_199;
      8'b11001000 : _zz_invSub_1 = invSboxRom_200;
      8'b11001001 : _zz_invSub_1 = invSboxRom_201;
      8'b11001010 : _zz_invSub_1 = invSboxRom_202;
      8'b11001011 : _zz_invSub_1 = invSboxRom_203;
      8'b11001100 : _zz_invSub_1 = invSboxRom_204;
      8'b11001101 : _zz_invSub_1 = invSboxRom_205;
      8'b11001110 : _zz_invSub_1 = invSboxRom_206;
      8'b11001111 : _zz_invSub_1 = invSboxRom_207;
      8'b11010000 : _zz_invSub_1 = invSboxRom_208;
      8'b11010001 : _zz_invSub_1 = invSboxRom_209;
      8'b11010010 : _zz_invSub_1 = invSboxRom_210;
      8'b11010011 : _zz_invSub_1 = invSboxRom_211;
      8'b11010100 : _zz_invSub_1 = invSboxRom_212;
      8'b11010101 : _zz_invSub_1 = invSboxRom_213;
      8'b11010110 : _zz_invSub_1 = invSboxRom_214;
      8'b11010111 : _zz_invSub_1 = invSboxRom_215;
      8'b11011000 : _zz_invSub_1 = invSboxRom_216;
      8'b11011001 : _zz_invSub_1 = invSboxRom_217;
      8'b11011010 : _zz_invSub_1 = invSboxRom_218;
      8'b11011011 : _zz_invSub_1 = invSboxRom_219;
      8'b11011100 : _zz_invSub_1 = invSboxRom_220;
      8'b11011101 : _zz_invSub_1 = invSboxRom_221;
      8'b11011110 : _zz_invSub_1 = invSboxRom_222;
      8'b11011111 : _zz_invSub_1 = invSboxRom_223;
      8'b11100000 : _zz_invSub_1 = invSboxRom_224;
      8'b11100001 : _zz_invSub_1 = invSboxRom_225;
      8'b11100010 : _zz_invSub_1 = invSboxRom_226;
      8'b11100011 : _zz_invSub_1 = invSboxRom_227;
      8'b11100100 : _zz_invSub_1 = invSboxRom_228;
      8'b11100101 : _zz_invSub_1 = invSboxRom_229;
      8'b11100110 : _zz_invSub_1 = invSboxRom_230;
      8'b11100111 : _zz_invSub_1 = invSboxRom_231;
      8'b11101000 : _zz_invSub_1 = invSboxRom_232;
      8'b11101001 : _zz_invSub_1 = invSboxRom_233;
      8'b11101010 : _zz_invSub_1 = invSboxRom_234;
      8'b11101011 : _zz_invSub_1 = invSboxRom_235;
      8'b11101100 : _zz_invSub_1 = invSboxRom_236;
      8'b11101101 : _zz_invSub_1 = invSboxRom_237;
      8'b11101110 : _zz_invSub_1 = invSboxRom_238;
      8'b11101111 : _zz_invSub_1 = invSboxRom_239;
      8'b11110000 : _zz_invSub_1 = invSboxRom_240;
      8'b11110001 : _zz_invSub_1 = invSboxRom_241;
      8'b11110010 : _zz_invSub_1 = invSboxRom_242;
      8'b11110011 : _zz_invSub_1 = invSboxRom_243;
      8'b11110100 : _zz_invSub_1 = invSboxRom_244;
      8'b11110101 : _zz_invSub_1 = invSboxRom_245;
      8'b11110110 : _zz_invSub_1 = invSboxRom_246;
      8'b11110111 : _zz_invSub_1 = invSboxRom_247;
      8'b11111000 : _zz_invSub_1 = invSboxRom_248;
      8'b11111001 : _zz_invSub_1 = invSboxRom_249;
      8'b11111010 : _zz_invSub_1 = invSboxRom_250;
      8'b11111011 : _zz_invSub_1 = invSboxRom_251;
      8'b11111100 : _zz_invSub_1 = invSboxRom_252;
      8'b11111101 : _zz_invSub_1 = invSboxRom_253;
      8'b11111110 : _zz_invSub_1 = invSboxRom_254;
      default : _zz_invSub_1 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_2)
      8'b00000000 : _zz_invSub_2 = invSboxRom_0;
      8'b00000001 : _zz_invSub_2 = invSboxRom_1;
      8'b00000010 : _zz_invSub_2 = invSboxRom_2;
      8'b00000011 : _zz_invSub_2 = invSboxRom_3;
      8'b00000100 : _zz_invSub_2 = invSboxRom_4;
      8'b00000101 : _zz_invSub_2 = invSboxRom_5;
      8'b00000110 : _zz_invSub_2 = invSboxRom_6;
      8'b00000111 : _zz_invSub_2 = invSboxRom_7;
      8'b00001000 : _zz_invSub_2 = invSboxRom_8;
      8'b00001001 : _zz_invSub_2 = invSboxRom_9;
      8'b00001010 : _zz_invSub_2 = invSboxRom_10;
      8'b00001011 : _zz_invSub_2 = invSboxRom_11;
      8'b00001100 : _zz_invSub_2 = invSboxRom_12;
      8'b00001101 : _zz_invSub_2 = invSboxRom_13;
      8'b00001110 : _zz_invSub_2 = invSboxRom_14;
      8'b00001111 : _zz_invSub_2 = invSboxRom_15;
      8'b00010000 : _zz_invSub_2 = invSboxRom_16;
      8'b00010001 : _zz_invSub_2 = invSboxRom_17;
      8'b00010010 : _zz_invSub_2 = invSboxRom_18;
      8'b00010011 : _zz_invSub_2 = invSboxRom_19;
      8'b00010100 : _zz_invSub_2 = invSboxRom_20;
      8'b00010101 : _zz_invSub_2 = invSboxRom_21;
      8'b00010110 : _zz_invSub_2 = invSboxRom_22;
      8'b00010111 : _zz_invSub_2 = invSboxRom_23;
      8'b00011000 : _zz_invSub_2 = invSboxRom_24;
      8'b00011001 : _zz_invSub_2 = invSboxRom_25;
      8'b00011010 : _zz_invSub_2 = invSboxRom_26;
      8'b00011011 : _zz_invSub_2 = invSboxRom_27;
      8'b00011100 : _zz_invSub_2 = invSboxRom_28;
      8'b00011101 : _zz_invSub_2 = invSboxRom_29;
      8'b00011110 : _zz_invSub_2 = invSboxRom_30;
      8'b00011111 : _zz_invSub_2 = invSboxRom_31;
      8'b00100000 : _zz_invSub_2 = invSboxRom_32;
      8'b00100001 : _zz_invSub_2 = invSboxRom_33;
      8'b00100010 : _zz_invSub_2 = invSboxRom_34;
      8'b00100011 : _zz_invSub_2 = invSboxRom_35;
      8'b00100100 : _zz_invSub_2 = invSboxRom_36;
      8'b00100101 : _zz_invSub_2 = invSboxRom_37;
      8'b00100110 : _zz_invSub_2 = invSboxRom_38;
      8'b00100111 : _zz_invSub_2 = invSboxRom_39;
      8'b00101000 : _zz_invSub_2 = invSboxRom_40;
      8'b00101001 : _zz_invSub_2 = invSboxRom_41;
      8'b00101010 : _zz_invSub_2 = invSboxRom_42;
      8'b00101011 : _zz_invSub_2 = invSboxRom_43;
      8'b00101100 : _zz_invSub_2 = invSboxRom_44;
      8'b00101101 : _zz_invSub_2 = invSboxRom_45;
      8'b00101110 : _zz_invSub_2 = invSboxRom_46;
      8'b00101111 : _zz_invSub_2 = invSboxRom_47;
      8'b00110000 : _zz_invSub_2 = invSboxRom_48;
      8'b00110001 : _zz_invSub_2 = invSboxRom_49;
      8'b00110010 : _zz_invSub_2 = invSboxRom_50;
      8'b00110011 : _zz_invSub_2 = invSboxRom_51;
      8'b00110100 : _zz_invSub_2 = invSboxRom_52;
      8'b00110101 : _zz_invSub_2 = invSboxRom_53;
      8'b00110110 : _zz_invSub_2 = invSboxRom_54;
      8'b00110111 : _zz_invSub_2 = invSboxRom_55;
      8'b00111000 : _zz_invSub_2 = invSboxRom_56;
      8'b00111001 : _zz_invSub_2 = invSboxRom_57;
      8'b00111010 : _zz_invSub_2 = invSboxRom_58;
      8'b00111011 : _zz_invSub_2 = invSboxRom_59;
      8'b00111100 : _zz_invSub_2 = invSboxRom_60;
      8'b00111101 : _zz_invSub_2 = invSboxRom_61;
      8'b00111110 : _zz_invSub_2 = invSboxRom_62;
      8'b00111111 : _zz_invSub_2 = invSboxRom_63;
      8'b01000000 : _zz_invSub_2 = invSboxRom_64;
      8'b01000001 : _zz_invSub_2 = invSboxRom_65;
      8'b01000010 : _zz_invSub_2 = invSboxRom_66;
      8'b01000011 : _zz_invSub_2 = invSboxRom_67;
      8'b01000100 : _zz_invSub_2 = invSboxRom_68;
      8'b01000101 : _zz_invSub_2 = invSboxRom_69;
      8'b01000110 : _zz_invSub_2 = invSboxRom_70;
      8'b01000111 : _zz_invSub_2 = invSboxRom_71;
      8'b01001000 : _zz_invSub_2 = invSboxRom_72;
      8'b01001001 : _zz_invSub_2 = invSboxRom_73;
      8'b01001010 : _zz_invSub_2 = invSboxRom_74;
      8'b01001011 : _zz_invSub_2 = invSboxRom_75;
      8'b01001100 : _zz_invSub_2 = invSboxRom_76;
      8'b01001101 : _zz_invSub_2 = invSboxRom_77;
      8'b01001110 : _zz_invSub_2 = invSboxRom_78;
      8'b01001111 : _zz_invSub_2 = invSboxRom_79;
      8'b01010000 : _zz_invSub_2 = invSboxRom_80;
      8'b01010001 : _zz_invSub_2 = invSboxRom_81;
      8'b01010010 : _zz_invSub_2 = invSboxRom_82;
      8'b01010011 : _zz_invSub_2 = invSboxRom_83;
      8'b01010100 : _zz_invSub_2 = invSboxRom_84;
      8'b01010101 : _zz_invSub_2 = invSboxRom_85;
      8'b01010110 : _zz_invSub_2 = invSboxRom_86;
      8'b01010111 : _zz_invSub_2 = invSboxRom_87;
      8'b01011000 : _zz_invSub_2 = invSboxRom_88;
      8'b01011001 : _zz_invSub_2 = invSboxRom_89;
      8'b01011010 : _zz_invSub_2 = invSboxRom_90;
      8'b01011011 : _zz_invSub_2 = invSboxRom_91;
      8'b01011100 : _zz_invSub_2 = invSboxRom_92;
      8'b01011101 : _zz_invSub_2 = invSboxRom_93;
      8'b01011110 : _zz_invSub_2 = invSboxRom_94;
      8'b01011111 : _zz_invSub_2 = invSboxRom_95;
      8'b01100000 : _zz_invSub_2 = invSboxRom_96;
      8'b01100001 : _zz_invSub_2 = invSboxRom_97;
      8'b01100010 : _zz_invSub_2 = invSboxRom_98;
      8'b01100011 : _zz_invSub_2 = invSboxRom_99;
      8'b01100100 : _zz_invSub_2 = invSboxRom_100;
      8'b01100101 : _zz_invSub_2 = invSboxRom_101;
      8'b01100110 : _zz_invSub_2 = invSboxRom_102;
      8'b01100111 : _zz_invSub_2 = invSboxRom_103;
      8'b01101000 : _zz_invSub_2 = invSboxRom_104;
      8'b01101001 : _zz_invSub_2 = invSboxRom_105;
      8'b01101010 : _zz_invSub_2 = invSboxRom_106;
      8'b01101011 : _zz_invSub_2 = invSboxRom_107;
      8'b01101100 : _zz_invSub_2 = invSboxRom_108;
      8'b01101101 : _zz_invSub_2 = invSboxRom_109;
      8'b01101110 : _zz_invSub_2 = invSboxRom_110;
      8'b01101111 : _zz_invSub_2 = invSboxRom_111;
      8'b01110000 : _zz_invSub_2 = invSboxRom_112;
      8'b01110001 : _zz_invSub_2 = invSboxRom_113;
      8'b01110010 : _zz_invSub_2 = invSboxRom_114;
      8'b01110011 : _zz_invSub_2 = invSboxRom_115;
      8'b01110100 : _zz_invSub_2 = invSboxRom_116;
      8'b01110101 : _zz_invSub_2 = invSboxRom_117;
      8'b01110110 : _zz_invSub_2 = invSboxRom_118;
      8'b01110111 : _zz_invSub_2 = invSboxRom_119;
      8'b01111000 : _zz_invSub_2 = invSboxRom_120;
      8'b01111001 : _zz_invSub_2 = invSboxRom_121;
      8'b01111010 : _zz_invSub_2 = invSboxRom_122;
      8'b01111011 : _zz_invSub_2 = invSboxRom_123;
      8'b01111100 : _zz_invSub_2 = invSboxRom_124;
      8'b01111101 : _zz_invSub_2 = invSboxRom_125;
      8'b01111110 : _zz_invSub_2 = invSboxRom_126;
      8'b01111111 : _zz_invSub_2 = invSboxRom_127;
      8'b10000000 : _zz_invSub_2 = invSboxRom_128;
      8'b10000001 : _zz_invSub_2 = invSboxRom_129;
      8'b10000010 : _zz_invSub_2 = invSboxRom_130;
      8'b10000011 : _zz_invSub_2 = invSboxRom_131;
      8'b10000100 : _zz_invSub_2 = invSboxRom_132;
      8'b10000101 : _zz_invSub_2 = invSboxRom_133;
      8'b10000110 : _zz_invSub_2 = invSboxRom_134;
      8'b10000111 : _zz_invSub_2 = invSboxRom_135;
      8'b10001000 : _zz_invSub_2 = invSboxRom_136;
      8'b10001001 : _zz_invSub_2 = invSboxRom_137;
      8'b10001010 : _zz_invSub_2 = invSboxRom_138;
      8'b10001011 : _zz_invSub_2 = invSboxRom_139;
      8'b10001100 : _zz_invSub_2 = invSboxRom_140;
      8'b10001101 : _zz_invSub_2 = invSboxRom_141;
      8'b10001110 : _zz_invSub_2 = invSboxRom_142;
      8'b10001111 : _zz_invSub_2 = invSboxRom_143;
      8'b10010000 : _zz_invSub_2 = invSboxRom_144;
      8'b10010001 : _zz_invSub_2 = invSboxRom_145;
      8'b10010010 : _zz_invSub_2 = invSboxRom_146;
      8'b10010011 : _zz_invSub_2 = invSboxRom_147;
      8'b10010100 : _zz_invSub_2 = invSboxRom_148;
      8'b10010101 : _zz_invSub_2 = invSboxRom_149;
      8'b10010110 : _zz_invSub_2 = invSboxRom_150;
      8'b10010111 : _zz_invSub_2 = invSboxRom_151;
      8'b10011000 : _zz_invSub_2 = invSboxRom_152;
      8'b10011001 : _zz_invSub_2 = invSboxRom_153;
      8'b10011010 : _zz_invSub_2 = invSboxRom_154;
      8'b10011011 : _zz_invSub_2 = invSboxRom_155;
      8'b10011100 : _zz_invSub_2 = invSboxRom_156;
      8'b10011101 : _zz_invSub_2 = invSboxRom_157;
      8'b10011110 : _zz_invSub_2 = invSboxRom_158;
      8'b10011111 : _zz_invSub_2 = invSboxRom_159;
      8'b10100000 : _zz_invSub_2 = invSboxRom_160;
      8'b10100001 : _zz_invSub_2 = invSboxRom_161;
      8'b10100010 : _zz_invSub_2 = invSboxRom_162;
      8'b10100011 : _zz_invSub_2 = invSboxRom_163;
      8'b10100100 : _zz_invSub_2 = invSboxRom_164;
      8'b10100101 : _zz_invSub_2 = invSboxRom_165;
      8'b10100110 : _zz_invSub_2 = invSboxRom_166;
      8'b10100111 : _zz_invSub_2 = invSboxRom_167;
      8'b10101000 : _zz_invSub_2 = invSboxRom_168;
      8'b10101001 : _zz_invSub_2 = invSboxRom_169;
      8'b10101010 : _zz_invSub_2 = invSboxRom_170;
      8'b10101011 : _zz_invSub_2 = invSboxRom_171;
      8'b10101100 : _zz_invSub_2 = invSboxRom_172;
      8'b10101101 : _zz_invSub_2 = invSboxRom_173;
      8'b10101110 : _zz_invSub_2 = invSboxRom_174;
      8'b10101111 : _zz_invSub_2 = invSboxRom_175;
      8'b10110000 : _zz_invSub_2 = invSboxRom_176;
      8'b10110001 : _zz_invSub_2 = invSboxRom_177;
      8'b10110010 : _zz_invSub_2 = invSboxRom_178;
      8'b10110011 : _zz_invSub_2 = invSboxRom_179;
      8'b10110100 : _zz_invSub_2 = invSboxRom_180;
      8'b10110101 : _zz_invSub_2 = invSboxRom_181;
      8'b10110110 : _zz_invSub_2 = invSboxRom_182;
      8'b10110111 : _zz_invSub_2 = invSboxRom_183;
      8'b10111000 : _zz_invSub_2 = invSboxRom_184;
      8'b10111001 : _zz_invSub_2 = invSboxRom_185;
      8'b10111010 : _zz_invSub_2 = invSboxRom_186;
      8'b10111011 : _zz_invSub_2 = invSboxRom_187;
      8'b10111100 : _zz_invSub_2 = invSboxRom_188;
      8'b10111101 : _zz_invSub_2 = invSboxRom_189;
      8'b10111110 : _zz_invSub_2 = invSboxRom_190;
      8'b10111111 : _zz_invSub_2 = invSboxRom_191;
      8'b11000000 : _zz_invSub_2 = invSboxRom_192;
      8'b11000001 : _zz_invSub_2 = invSboxRom_193;
      8'b11000010 : _zz_invSub_2 = invSboxRom_194;
      8'b11000011 : _zz_invSub_2 = invSboxRom_195;
      8'b11000100 : _zz_invSub_2 = invSboxRom_196;
      8'b11000101 : _zz_invSub_2 = invSboxRom_197;
      8'b11000110 : _zz_invSub_2 = invSboxRom_198;
      8'b11000111 : _zz_invSub_2 = invSboxRom_199;
      8'b11001000 : _zz_invSub_2 = invSboxRom_200;
      8'b11001001 : _zz_invSub_2 = invSboxRom_201;
      8'b11001010 : _zz_invSub_2 = invSboxRom_202;
      8'b11001011 : _zz_invSub_2 = invSboxRom_203;
      8'b11001100 : _zz_invSub_2 = invSboxRom_204;
      8'b11001101 : _zz_invSub_2 = invSboxRom_205;
      8'b11001110 : _zz_invSub_2 = invSboxRom_206;
      8'b11001111 : _zz_invSub_2 = invSboxRom_207;
      8'b11010000 : _zz_invSub_2 = invSboxRom_208;
      8'b11010001 : _zz_invSub_2 = invSboxRom_209;
      8'b11010010 : _zz_invSub_2 = invSboxRom_210;
      8'b11010011 : _zz_invSub_2 = invSboxRom_211;
      8'b11010100 : _zz_invSub_2 = invSboxRom_212;
      8'b11010101 : _zz_invSub_2 = invSboxRom_213;
      8'b11010110 : _zz_invSub_2 = invSboxRom_214;
      8'b11010111 : _zz_invSub_2 = invSboxRom_215;
      8'b11011000 : _zz_invSub_2 = invSboxRom_216;
      8'b11011001 : _zz_invSub_2 = invSboxRom_217;
      8'b11011010 : _zz_invSub_2 = invSboxRom_218;
      8'b11011011 : _zz_invSub_2 = invSboxRom_219;
      8'b11011100 : _zz_invSub_2 = invSboxRom_220;
      8'b11011101 : _zz_invSub_2 = invSboxRom_221;
      8'b11011110 : _zz_invSub_2 = invSboxRom_222;
      8'b11011111 : _zz_invSub_2 = invSboxRom_223;
      8'b11100000 : _zz_invSub_2 = invSboxRom_224;
      8'b11100001 : _zz_invSub_2 = invSboxRom_225;
      8'b11100010 : _zz_invSub_2 = invSboxRom_226;
      8'b11100011 : _zz_invSub_2 = invSboxRom_227;
      8'b11100100 : _zz_invSub_2 = invSboxRom_228;
      8'b11100101 : _zz_invSub_2 = invSboxRom_229;
      8'b11100110 : _zz_invSub_2 = invSboxRom_230;
      8'b11100111 : _zz_invSub_2 = invSboxRom_231;
      8'b11101000 : _zz_invSub_2 = invSboxRom_232;
      8'b11101001 : _zz_invSub_2 = invSboxRom_233;
      8'b11101010 : _zz_invSub_2 = invSboxRom_234;
      8'b11101011 : _zz_invSub_2 = invSboxRom_235;
      8'b11101100 : _zz_invSub_2 = invSboxRom_236;
      8'b11101101 : _zz_invSub_2 = invSboxRom_237;
      8'b11101110 : _zz_invSub_2 = invSboxRom_238;
      8'b11101111 : _zz_invSub_2 = invSboxRom_239;
      8'b11110000 : _zz_invSub_2 = invSboxRom_240;
      8'b11110001 : _zz_invSub_2 = invSboxRom_241;
      8'b11110010 : _zz_invSub_2 = invSboxRom_242;
      8'b11110011 : _zz_invSub_2 = invSboxRom_243;
      8'b11110100 : _zz_invSub_2 = invSboxRom_244;
      8'b11110101 : _zz_invSub_2 = invSboxRom_245;
      8'b11110110 : _zz_invSub_2 = invSboxRom_246;
      8'b11110111 : _zz_invSub_2 = invSboxRom_247;
      8'b11111000 : _zz_invSub_2 = invSboxRom_248;
      8'b11111001 : _zz_invSub_2 = invSboxRom_249;
      8'b11111010 : _zz_invSub_2 = invSboxRom_250;
      8'b11111011 : _zz_invSub_2 = invSboxRom_251;
      8'b11111100 : _zz_invSub_2 = invSboxRom_252;
      8'b11111101 : _zz_invSub_2 = invSboxRom_253;
      8'b11111110 : _zz_invSub_2 = invSboxRom_254;
      default : _zz_invSub_2 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_3)
      8'b00000000 : _zz_invSub_3 = invSboxRom_0;
      8'b00000001 : _zz_invSub_3 = invSboxRom_1;
      8'b00000010 : _zz_invSub_3 = invSboxRom_2;
      8'b00000011 : _zz_invSub_3 = invSboxRom_3;
      8'b00000100 : _zz_invSub_3 = invSboxRom_4;
      8'b00000101 : _zz_invSub_3 = invSboxRom_5;
      8'b00000110 : _zz_invSub_3 = invSboxRom_6;
      8'b00000111 : _zz_invSub_3 = invSboxRom_7;
      8'b00001000 : _zz_invSub_3 = invSboxRom_8;
      8'b00001001 : _zz_invSub_3 = invSboxRom_9;
      8'b00001010 : _zz_invSub_3 = invSboxRom_10;
      8'b00001011 : _zz_invSub_3 = invSboxRom_11;
      8'b00001100 : _zz_invSub_3 = invSboxRom_12;
      8'b00001101 : _zz_invSub_3 = invSboxRom_13;
      8'b00001110 : _zz_invSub_3 = invSboxRom_14;
      8'b00001111 : _zz_invSub_3 = invSboxRom_15;
      8'b00010000 : _zz_invSub_3 = invSboxRom_16;
      8'b00010001 : _zz_invSub_3 = invSboxRom_17;
      8'b00010010 : _zz_invSub_3 = invSboxRom_18;
      8'b00010011 : _zz_invSub_3 = invSboxRom_19;
      8'b00010100 : _zz_invSub_3 = invSboxRom_20;
      8'b00010101 : _zz_invSub_3 = invSboxRom_21;
      8'b00010110 : _zz_invSub_3 = invSboxRom_22;
      8'b00010111 : _zz_invSub_3 = invSboxRom_23;
      8'b00011000 : _zz_invSub_3 = invSboxRom_24;
      8'b00011001 : _zz_invSub_3 = invSboxRom_25;
      8'b00011010 : _zz_invSub_3 = invSboxRom_26;
      8'b00011011 : _zz_invSub_3 = invSboxRom_27;
      8'b00011100 : _zz_invSub_3 = invSboxRom_28;
      8'b00011101 : _zz_invSub_3 = invSboxRom_29;
      8'b00011110 : _zz_invSub_3 = invSboxRom_30;
      8'b00011111 : _zz_invSub_3 = invSboxRom_31;
      8'b00100000 : _zz_invSub_3 = invSboxRom_32;
      8'b00100001 : _zz_invSub_3 = invSboxRom_33;
      8'b00100010 : _zz_invSub_3 = invSboxRom_34;
      8'b00100011 : _zz_invSub_3 = invSboxRom_35;
      8'b00100100 : _zz_invSub_3 = invSboxRom_36;
      8'b00100101 : _zz_invSub_3 = invSboxRom_37;
      8'b00100110 : _zz_invSub_3 = invSboxRom_38;
      8'b00100111 : _zz_invSub_3 = invSboxRom_39;
      8'b00101000 : _zz_invSub_3 = invSboxRom_40;
      8'b00101001 : _zz_invSub_3 = invSboxRom_41;
      8'b00101010 : _zz_invSub_3 = invSboxRom_42;
      8'b00101011 : _zz_invSub_3 = invSboxRom_43;
      8'b00101100 : _zz_invSub_3 = invSboxRom_44;
      8'b00101101 : _zz_invSub_3 = invSboxRom_45;
      8'b00101110 : _zz_invSub_3 = invSboxRom_46;
      8'b00101111 : _zz_invSub_3 = invSboxRom_47;
      8'b00110000 : _zz_invSub_3 = invSboxRom_48;
      8'b00110001 : _zz_invSub_3 = invSboxRom_49;
      8'b00110010 : _zz_invSub_3 = invSboxRom_50;
      8'b00110011 : _zz_invSub_3 = invSboxRom_51;
      8'b00110100 : _zz_invSub_3 = invSboxRom_52;
      8'b00110101 : _zz_invSub_3 = invSboxRom_53;
      8'b00110110 : _zz_invSub_3 = invSboxRom_54;
      8'b00110111 : _zz_invSub_3 = invSboxRom_55;
      8'b00111000 : _zz_invSub_3 = invSboxRom_56;
      8'b00111001 : _zz_invSub_3 = invSboxRom_57;
      8'b00111010 : _zz_invSub_3 = invSboxRom_58;
      8'b00111011 : _zz_invSub_3 = invSboxRom_59;
      8'b00111100 : _zz_invSub_3 = invSboxRom_60;
      8'b00111101 : _zz_invSub_3 = invSboxRom_61;
      8'b00111110 : _zz_invSub_3 = invSboxRom_62;
      8'b00111111 : _zz_invSub_3 = invSboxRom_63;
      8'b01000000 : _zz_invSub_3 = invSboxRom_64;
      8'b01000001 : _zz_invSub_3 = invSboxRom_65;
      8'b01000010 : _zz_invSub_3 = invSboxRom_66;
      8'b01000011 : _zz_invSub_3 = invSboxRom_67;
      8'b01000100 : _zz_invSub_3 = invSboxRom_68;
      8'b01000101 : _zz_invSub_3 = invSboxRom_69;
      8'b01000110 : _zz_invSub_3 = invSboxRom_70;
      8'b01000111 : _zz_invSub_3 = invSboxRom_71;
      8'b01001000 : _zz_invSub_3 = invSboxRom_72;
      8'b01001001 : _zz_invSub_3 = invSboxRom_73;
      8'b01001010 : _zz_invSub_3 = invSboxRom_74;
      8'b01001011 : _zz_invSub_3 = invSboxRom_75;
      8'b01001100 : _zz_invSub_3 = invSboxRom_76;
      8'b01001101 : _zz_invSub_3 = invSboxRom_77;
      8'b01001110 : _zz_invSub_3 = invSboxRom_78;
      8'b01001111 : _zz_invSub_3 = invSboxRom_79;
      8'b01010000 : _zz_invSub_3 = invSboxRom_80;
      8'b01010001 : _zz_invSub_3 = invSboxRom_81;
      8'b01010010 : _zz_invSub_3 = invSboxRom_82;
      8'b01010011 : _zz_invSub_3 = invSboxRom_83;
      8'b01010100 : _zz_invSub_3 = invSboxRom_84;
      8'b01010101 : _zz_invSub_3 = invSboxRom_85;
      8'b01010110 : _zz_invSub_3 = invSboxRom_86;
      8'b01010111 : _zz_invSub_3 = invSboxRom_87;
      8'b01011000 : _zz_invSub_3 = invSboxRom_88;
      8'b01011001 : _zz_invSub_3 = invSboxRom_89;
      8'b01011010 : _zz_invSub_3 = invSboxRom_90;
      8'b01011011 : _zz_invSub_3 = invSboxRom_91;
      8'b01011100 : _zz_invSub_3 = invSboxRom_92;
      8'b01011101 : _zz_invSub_3 = invSboxRom_93;
      8'b01011110 : _zz_invSub_3 = invSboxRom_94;
      8'b01011111 : _zz_invSub_3 = invSboxRom_95;
      8'b01100000 : _zz_invSub_3 = invSboxRom_96;
      8'b01100001 : _zz_invSub_3 = invSboxRom_97;
      8'b01100010 : _zz_invSub_3 = invSboxRom_98;
      8'b01100011 : _zz_invSub_3 = invSboxRom_99;
      8'b01100100 : _zz_invSub_3 = invSboxRom_100;
      8'b01100101 : _zz_invSub_3 = invSboxRom_101;
      8'b01100110 : _zz_invSub_3 = invSboxRom_102;
      8'b01100111 : _zz_invSub_3 = invSboxRom_103;
      8'b01101000 : _zz_invSub_3 = invSboxRom_104;
      8'b01101001 : _zz_invSub_3 = invSboxRom_105;
      8'b01101010 : _zz_invSub_3 = invSboxRom_106;
      8'b01101011 : _zz_invSub_3 = invSboxRom_107;
      8'b01101100 : _zz_invSub_3 = invSboxRom_108;
      8'b01101101 : _zz_invSub_3 = invSboxRom_109;
      8'b01101110 : _zz_invSub_3 = invSboxRom_110;
      8'b01101111 : _zz_invSub_3 = invSboxRom_111;
      8'b01110000 : _zz_invSub_3 = invSboxRom_112;
      8'b01110001 : _zz_invSub_3 = invSboxRom_113;
      8'b01110010 : _zz_invSub_3 = invSboxRom_114;
      8'b01110011 : _zz_invSub_3 = invSboxRom_115;
      8'b01110100 : _zz_invSub_3 = invSboxRom_116;
      8'b01110101 : _zz_invSub_3 = invSboxRom_117;
      8'b01110110 : _zz_invSub_3 = invSboxRom_118;
      8'b01110111 : _zz_invSub_3 = invSboxRom_119;
      8'b01111000 : _zz_invSub_3 = invSboxRom_120;
      8'b01111001 : _zz_invSub_3 = invSboxRom_121;
      8'b01111010 : _zz_invSub_3 = invSboxRom_122;
      8'b01111011 : _zz_invSub_3 = invSboxRom_123;
      8'b01111100 : _zz_invSub_3 = invSboxRom_124;
      8'b01111101 : _zz_invSub_3 = invSboxRom_125;
      8'b01111110 : _zz_invSub_3 = invSboxRom_126;
      8'b01111111 : _zz_invSub_3 = invSboxRom_127;
      8'b10000000 : _zz_invSub_3 = invSboxRom_128;
      8'b10000001 : _zz_invSub_3 = invSboxRom_129;
      8'b10000010 : _zz_invSub_3 = invSboxRom_130;
      8'b10000011 : _zz_invSub_3 = invSboxRom_131;
      8'b10000100 : _zz_invSub_3 = invSboxRom_132;
      8'b10000101 : _zz_invSub_3 = invSboxRom_133;
      8'b10000110 : _zz_invSub_3 = invSboxRom_134;
      8'b10000111 : _zz_invSub_3 = invSboxRom_135;
      8'b10001000 : _zz_invSub_3 = invSboxRom_136;
      8'b10001001 : _zz_invSub_3 = invSboxRom_137;
      8'b10001010 : _zz_invSub_3 = invSboxRom_138;
      8'b10001011 : _zz_invSub_3 = invSboxRom_139;
      8'b10001100 : _zz_invSub_3 = invSboxRom_140;
      8'b10001101 : _zz_invSub_3 = invSboxRom_141;
      8'b10001110 : _zz_invSub_3 = invSboxRom_142;
      8'b10001111 : _zz_invSub_3 = invSboxRom_143;
      8'b10010000 : _zz_invSub_3 = invSboxRom_144;
      8'b10010001 : _zz_invSub_3 = invSboxRom_145;
      8'b10010010 : _zz_invSub_3 = invSboxRom_146;
      8'b10010011 : _zz_invSub_3 = invSboxRom_147;
      8'b10010100 : _zz_invSub_3 = invSboxRom_148;
      8'b10010101 : _zz_invSub_3 = invSboxRom_149;
      8'b10010110 : _zz_invSub_3 = invSboxRom_150;
      8'b10010111 : _zz_invSub_3 = invSboxRom_151;
      8'b10011000 : _zz_invSub_3 = invSboxRom_152;
      8'b10011001 : _zz_invSub_3 = invSboxRom_153;
      8'b10011010 : _zz_invSub_3 = invSboxRom_154;
      8'b10011011 : _zz_invSub_3 = invSboxRom_155;
      8'b10011100 : _zz_invSub_3 = invSboxRom_156;
      8'b10011101 : _zz_invSub_3 = invSboxRom_157;
      8'b10011110 : _zz_invSub_3 = invSboxRom_158;
      8'b10011111 : _zz_invSub_3 = invSboxRom_159;
      8'b10100000 : _zz_invSub_3 = invSboxRom_160;
      8'b10100001 : _zz_invSub_3 = invSboxRom_161;
      8'b10100010 : _zz_invSub_3 = invSboxRom_162;
      8'b10100011 : _zz_invSub_3 = invSboxRom_163;
      8'b10100100 : _zz_invSub_3 = invSboxRom_164;
      8'b10100101 : _zz_invSub_3 = invSboxRom_165;
      8'b10100110 : _zz_invSub_3 = invSboxRom_166;
      8'b10100111 : _zz_invSub_3 = invSboxRom_167;
      8'b10101000 : _zz_invSub_3 = invSboxRom_168;
      8'b10101001 : _zz_invSub_3 = invSboxRom_169;
      8'b10101010 : _zz_invSub_3 = invSboxRom_170;
      8'b10101011 : _zz_invSub_3 = invSboxRom_171;
      8'b10101100 : _zz_invSub_3 = invSboxRom_172;
      8'b10101101 : _zz_invSub_3 = invSboxRom_173;
      8'b10101110 : _zz_invSub_3 = invSboxRom_174;
      8'b10101111 : _zz_invSub_3 = invSboxRom_175;
      8'b10110000 : _zz_invSub_3 = invSboxRom_176;
      8'b10110001 : _zz_invSub_3 = invSboxRom_177;
      8'b10110010 : _zz_invSub_3 = invSboxRom_178;
      8'b10110011 : _zz_invSub_3 = invSboxRom_179;
      8'b10110100 : _zz_invSub_3 = invSboxRom_180;
      8'b10110101 : _zz_invSub_3 = invSboxRom_181;
      8'b10110110 : _zz_invSub_3 = invSboxRom_182;
      8'b10110111 : _zz_invSub_3 = invSboxRom_183;
      8'b10111000 : _zz_invSub_3 = invSboxRom_184;
      8'b10111001 : _zz_invSub_3 = invSboxRom_185;
      8'b10111010 : _zz_invSub_3 = invSboxRom_186;
      8'b10111011 : _zz_invSub_3 = invSboxRom_187;
      8'b10111100 : _zz_invSub_3 = invSboxRom_188;
      8'b10111101 : _zz_invSub_3 = invSboxRom_189;
      8'b10111110 : _zz_invSub_3 = invSboxRom_190;
      8'b10111111 : _zz_invSub_3 = invSboxRom_191;
      8'b11000000 : _zz_invSub_3 = invSboxRom_192;
      8'b11000001 : _zz_invSub_3 = invSboxRom_193;
      8'b11000010 : _zz_invSub_3 = invSboxRom_194;
      8'b11000011 : _zz_invSub_3 = invSboxRom_195;
      8'b11000100 : _zz_invSub_3 = invSboxRom_196;
      8'b11000101 : _zz_invSub_3 = invSboxRom_197;
      8'b11000110 : _zz_invSub_3 = invSboxRom_198;
      8'b11000111 : _zz_invSub_3 = invSboxRom_199;
      8'b11001000 : _zz_invSub_3 = invSboxRom_200;
      8'b11001001 : _zz_invSub_3 = invSboxRom_201;
      8'b11001010 : _zz_invSub_3 = invSboxRom_202;
      8'b11001011 : _zz_invSub_3 = invSboxRom_203;
      8'b11001100 : _zz_invSub_3 = invSboxRom_204;
      8'b11001101 : _zz_invSub_3 = invSboxRom_205;
      8'b11001110 : _zz_invSub_3 = invSboxRom_206;
      8'b11001111 : _zz_invSub_3 = invSboxRom_207;
      8'b11010000 : _zz_invSub_3 = invSboxRom_208;
      8'b11010001 : _zz_invSub_3 = invSboxRom_209;
      8'b11010010 : _zz_invSub_3 = invSboxRom_210;
      8'b11010011 : _zz_invSub_3 = invSboxRom_211;
      8'b11010100 : _zz_invSub_3 = invSboxRom_212;
      8'b11010101 : _zz_invSub_3 = invSboxRom_213;
      8'b11010110 : _zz_invSub_3 = invSboxRom_214;
      8'b11010111 : _zz_invSub_3 = invSboxRom_215;
      8'b11011000 : _zz_invSub_3 = invSboxRom_216;
      8'b11011001 : _zz_invSub_3 = invSboxRom_217;
      8'b11011010 : _zz_invSub_3 = invSboxRom_218;
      8'b11011011 : _zz_invSub_3 = invSboxRom_219;
      8'b11011100 : _zz_invSub_3 = invSboxRom_220;
      8'b11011101 : _zz_invSub_3 = invSboxRom_221;
      8'b11011110 : _zz_invSub_3 = invSboxRom_222;
      8'b11011111 : _zz_invSub_3 = invSboxRom_223;
      8'b11100000 : _zz_invSub_3 = invSboxRom_224;
      8'b11100001 : _zz_invSub_3 = invSboxRom_225;
      8'b11100010 : _zz_invSub_3 = invSboxRom_226;
      8'b11100011 : _zz_invSub_3 = invSboxRom_227;
      8'b11100100 : _zz_invSub_3 = invSboxRom_228;
      8'b11100101 : _zz_invSub_3 = invSboxRom_229;
      8'b11100110 : _zz_invSub_3 = invSboxRom_230;
      8'b11100111 : _zz_invSub_3 = invSboxRom_231;
      8'b11101000 : _zz_invSub_3 = invSboxRom_232;
      8'b11101001 : _zz_invSub_3 = invSboxRom_233;
      8'b11101010 : _zz_invSub_3 = invSboxRom_234;
      8'b11101011 : _zz_invSub_3 = invSboxRom_235;
      8'b11101100 : _zz_invSub_3 = invSboxRom_236;
      8'b11101101 : _zz_invSub_3 = invSboxRom_237;
      8'b11101110 : _zz_invSub_3 = invSboxRom_238;
      8'b11101111 : _zz_invSub_3 = invSboxRom_239;
      8'b11110000 : _zz_invSub_3 = invSboxRom_240;
      8'b11110001 : _zz_invSub_3 = invSboxRom_241;
      8'b11110010 : _zz_invSub_3 = invSboxRom_242;
      8'b11110011 : _zz_invSub_3 = invSboxRom_243;
      8'b11110100 : _zz_invSub_3 = invSboxRom_244;
      8'b11110101 : _zz_invSub_3 = invSboxRom_245;
      8'b11110110 : _zz_invSub_3 = invSboxRom_246;
      8'b11110111 : _zz_invSub_3 = invSboxRom_247;
      8'b11111000 : _zz_invSub_3 = invSboxRom_248;
      8'b11111001 : _zz_invSub_3 = invSboxRom_249;
      8'b11111010 : _zz_invSub_3 = invSboxRom_250;
      8'b11111011 : _zz_invSub_3 = invSboxRom_251;
      8'b11111100 : _zz_invSub_3 = invSboxRom_252;
      8'b11111101 : _zz_invSub_3 = invSboxRom_253;
      8'b11111110 : _zz_invSub_3 = invSboxRom_254;
      default : _zz_invSub_3 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_4)
      8'b00000000 : _zz_invSub_4 = invSboxRom_0;
      8'b00000001 : _zz_invSub_4 = invSboxRom_1;
      8'b00000010 : _zz_invSub_4 = invSboxRom_2;
      8'b00000011 : _zz_invSub_4 = invSboxRom_3;
      8'b00000100 : _zz_invSub_4 = invSboxRom_4;
      8'b00000101 : _zz_invSub_4 = invSboxRom_5;
      8'b00000110 : _zz_invSub_4 = invSboxRom_6;
      8'b00000111 : _zz_invSub_4 = invSboxRom_7;
      8'b00001000 : _zz_invSub_4 = invSboxRom_8;
      8'b00001001 : _zz_invSub_4 = invSboxRom_9;
      8'b00001010 : _zz_invSub_4 = invSboxRom_10;
      8'b00001011 : _zz_invSub_4 = invSboxRom_11;
      8'b00001100 : _zz_invSub_4 = invSboxRom_12;
      8'b00001101 : _zz_invSub_4 = invSboxRom_13;
      8'b00001110 : _zz_invSub_4 = invSboxRom_14;
      8'b00001111 : _zz_invSub_4 = invSboxRom_15;
      8'b00010000 : _zz_invSub_4 = invSboxRom_16;
      8'b00010001 : _zz_invSub_4 = invSboxRom_17;
      8'b00010010 : _zz_invSub_4 = invSboxRom_18;
      8'b00010011 : _zz_invSub_4 = invSboxRom_19;
      8'b00010100 : _zz_invSub_4 = invSboxRom_20;
      8'b00010101 : _zz_invSub_4 = invSboxRom_21;
      8'b00010110 : _zz_invSub_4 = invSboxRom_22;
      8'b00010111 : _zz_invSub_4 = invSboxRom_23;
      8'b00011000 : _zz_invSub_4 = invSboxRom_24;
      8'b00011001 : _zz_invSub_4 = invSboxRom_25;
      8'b00011010 : _zz_invSub_4 = invSboxRom_26;
      8'b00011011 : _zz_invSub_4 = invSboxRom_27;
      8'b00011100 : _zz_invSub_4 = invSboxRom_28;
      8'b00011101 : _zz_invSub_4 = invSboxRom_29;
      8'b00011110 : _zz_invSub_4 = invSboxRom_30;
      8'b00011111 : _zz_invSub_4 = invSboxRom_31;
      8'b00100000 : _zz_invSub_4 = invSboxRom_32;
      8'b00100001 : _zz_invSub_4 = invSboxRom_33;
      8'b00100010 : _zz_invSub_4 = invSboxRom_34;
      8'b00100011 : _zz_invSub_4 = invSboxRom_35;
      8'b00100100 : _zz_invSub_4 = invSboxRom_36;
      8'b00100101 : _zz_invSub_4 = invSboxRom_37;
      8'b00100110 : _zz_invSub_4 = invSboxRom_38;
      8'b00100111 : _zz_invSub_4 = invSboxRom_39;
      8'b00101000 : _zz_invSub_4 = invSboxRom_40;
      8'b00101001 : _zz_invSub_4 = invSboxRom_41;
      8'b00101010 : _zz_invSub_4 = invSboxRom_42;
      8'b00101011 : _zz_invSub_4 = invSboxRom_43;
      8'b00101100 : _zz_invSub_4 = invSboxRom_44;
      8'b00101101 : _zz_invSub_4 = invSboxRom_45;
      8'b00101110 : _zz_invSub_4 = invSboxRom_46;
      8'b00101111 : _zz_invSub_4 = invSboxRom_47;
      8'b00110000 : _zz_invSub_4 = invSboxRom_48;
      8'b00110001 : _zz_invSub_4 = invSboxRom_49;
      8'b00110010 : _zz_invSub_4 = invSboxRom_50;
      8'b00110011 : _zz_invSub_4 = invSboxRom_51;
      8'b00110100 : _zz_invSub_4 = invSboxRom_52;
      8'b00110101 : _zz_invSub_4 = invSboxRom_53;
      8'b00110110 : _zz_invSub_4 = invSboxRom_54;
      8'b00110111 : _zz_invSub_4 = invSboxRom_55;
      8'b00111000 : _zz_invSub_4 = invSboxRom_56;
      8'b00111001 : _zz_invSub_4 = invSboxRom_57;
      8'b00111010 : _zz_invSub_4 = invSboxRom_58;
      8'b00111011 : _zz_invSub_4 = invSboxRom_59;
      8'b00111100 : _zz_invSub_4 = invSboxRom_60;
      8'b00111101 : _zz_invSub_4 = invSboxRom_61;
      8'b00111110 : _zz_invSub_4 = invSboxRom_62;
      8'b00111111 : _zz_invSub_4 = invSboxRom_63;
      8'b01000000 : _zz_invSub_4 = invSboxRom_64;
      8'b01000001 : _zz_invSub_4 = invSboxRom_65;
      8'b01000010 : _zz_invSub_4 = invSboxRom_66;
      8'b01000011 : _zz_invSub_4 = invSboxRom_67;
      8'b01000100 : _zz_invSub_4 = invSboxRom_68;
      8'b01000101 : _zz_invSub_4 = invSboxRom_69;
      8'b01000110 : _zz_invSub_4 = invSboxRom_70;
      8'b01000111 : _zz_invSub_4 = invSboxRom_71;
      8'b01001000 : _zz_invSub_4 = invSboxRom_72;
      8'b01001001 : _zz_invSub_4 = invSboxRom_73;
      8'b01001010 : _zz_invSub_4 = invSboxRom_74;
      8'b01001011 : _zz_invSub_4 = invSboxRom_75;
      8'b01001100 : _zz_invSub_4 = invSboxRom_76;
      8'b01001101 : _zz_invSub_4 = invSboxRom_77;
      8'b01001110 : _zz_invSub_4 = invSboxRom_78;
      8'b01001111 : _zz_invSub_4 = invSboxRom_79;
      8'b01010000 : _zz_invSub_4 = invSboxRom_80;
      8'b01010001 : _zz_invSub_4 = invSboxRom_81;
      8'b01010010 : _zz_invSub_4 = invSboxRom_82;
      8'b01010011 : _zz_invSub_4 = invSboxRom_83;
      8'b01010100 : _zz_invSub_4 = invSboxRom_84;
      8'b01010101 : _zz_invSub_4 = invSboxRom_85;
      8'b01010110 : _zz_invSub_4 = invSboxRom_86;
      8'b01010111 : _zz_invSub_4 = invSboxRom_87;
      8'b01011000 : _zz_invSub_4 = invSboxRom_88;
      8'b01011001 : _zz_invSub_4 = invSboxRom_89;
      8'b01011010 : _zz_invSub_4 = invSboxRom_90;
      8'b01011011 : _zz_invSub_4 = invSboxRom_91;
      8'b01011100 : _zz_invSub_4 = invSboxRom_92;
      8'b01011101 : _zz_invSub_4 = invSboxRom_93;
      8'b01011110 : _zz_invSub_4 = invSboxRom_94;
      8'b01011111 : _zz_invSub_4 = invSboxRom_95;
      8'b01100000 : _zz_invSub_4 = invSboxRom_96;
      8'b01100001 : _zz_invSub_4 = invSboxRom_97;
      8'b01100010 : _zz_invSub_4 = invSboxRom_98;
      8'b01100011 : _zz_invSub_4 = invSboxRom_99;
      8'b01100100 : _zz_invSub_4 = invSboxRom_100;
      8'b01100101 : _zz_invSub_4 = invSboxRom_101;
      8'b01100110 : _zz_invSub_4 = invSboxRom_102;
      8'b01100111 : _zz_invSub_4 = invSboxRom_103;
      8'b01101000 : _zz_invSub_4 = invSboxRom_104;
      8'b01101001 : _zz_invSub_4 = invSboxRom_105;
      8'b01101010 : _zz_invSub_4 = invSboxRom_106;
      8'b01101011 : _zz_invSub_4 = invSboxRom_107;
      8'b01101100 : _zz_invSub_4 = invSboxRom_108;
      8'b01101101 : _zz_invSub_4 = invSboxRom_109;
      8'b01101110 : _zz_invSub_4 = invSboxRom_110;
      8'b01101111 : _zz_invSub_4 = invSboxRom_111;
      8'b01110000 : _zz_invSub_4 = invSboxRom_112;
      8'b01110001 : _zz_invSub_4 = invSboxRom_113;
      8'b01110010 : _zz_invSub_4 = invSboxRom_114;
      8'b01110011 : _zz_invSub_4 = invSboxRom_115;
      8'b01110100 : _zz_invSub_4 = invSboxRom_116;
      8'b01110101 : _zz_invSub_4 = invSboxRom_117;
      8'b01110110 : _zz_invSub_4 = invSboxRom_118;
      8'b01110111 : _zz_invSub_4 = invSboxRom_119;
      8'b01111000 : _zz_invSub_4 = invSboxRom_120;
      8'b01111001 : _zz_invSub_4 = invSboxRom_121;
      8'b01111010 : _zz_invSub_4 = invSboxRom_122;
      8'b01111011 : _zz_invSub_4 = invSboxRom_123;
      8'b01111100 : _zz_invSub_4 = invSboxRom_124;
      8'b01111101 : _zz_invSub_4 = invSboxRom_125;
      8'b01111110 : _zz_invSub_4 = invSboxRom_126;
      8'b01111111 : _zz_invSub_4 = invSboxRom_127;
      8'b10000000 : _zz_invSub_4 = invSboxRom_128;
      8'b10000001 : _zz_invSub_4 = invSboxRom_129;
      8'b10000010 : _zz_invSub_4 = invSboxRom_130;
      8'b10000011 : _zz_invSub_4 = invSboxRom_131;
      8'b10000100 : _zz_invSub_4 = invSboxRom_132;
      8'b10000101 : _zz_invSub_4 = invSboxRom_133;
      8'b10000110 : _zz_invSub_4 = invSboxRom_134;
      8'b10000111 : _zz_invSub_4 = invSboxRom_135;
      8'b10001000 : _zz_invSub_4 = invSboxRom_136;
      8'b10001001 : _zz_invSub_4 = invSboxRom_137;
      8'b10001010 : _zz_invSub_4 = invSboxRom_138;
      8'b10001011 : _zz_invSub_4 = invSboxRom_139;
      8'b10001100 : _zz_invSub_4 = invSboxRom_140;
      8'b10001101 : _zz_invSub_4 = invSboxRom_141;
      8'b10001110 : _zz_invSub_4 = invSboxRom_142;
      8'b10001111 : _zz_invSub_4 = invSboxRom_143;
      8'b10010000 : _zz_invSub_4 = invSboxRom_144;
      8'b10010001 : _zz_invSub_4 = invSboxRom_145;
      8'b10010010 : _zz_invSub_4 = invSboxRom_146;
      8'b10010011 : _zz_invSub_4 = invSboxRom_147;
      8'b10010100 : _zz_invSub_4 = invSboxRom_148;
      8'b10010101 : _zz_invSub_4 = invSboxRom_149;
      8'b10010110 : _zz_invSub_4 = invSboxRom_150;
      8'b10010111 : _zz_invSub_4 = invSboxRom_151;
      8'b10011000 : _zz_invSub_4 = invSboxRom_152;
      8'b10011001 : _zz_invSub_4 = invSboxRom_153;
      8'b10011010 : _zz_invSub_4 = invSboxRom_154;
      8'b10011011 : _zz_invSub_4 = invSboxRom_155;
      8'b10011100 : _zz_invSub_4 = invSboxRom_156;
      8'b10011101 : _zz_invSub_4 = invSboxRom_157;
      8'b10011110 : _zz_invSub_4 = invSboxRom_158;
      8'b10011111 : _zz_invSub_4 = invSboxRom_159;
      8'b10100000 : _zz_invSub_4 = invSboxRom_160;
      8'b10100001 : _zz_invSub_4 = invSboxRom_161;
      8'b10100010 : _zz_invSub_4 = invSboxRom_162;
      8'b10100011 : _zz_invSub_4 = invSboxRom_163;
      8'b10100100 : _zz_invSub_4 = invSboxRom_164;
      8'b10100101 : _zz_invSub_4 = invSboxRom_165;
      8'b10100110 : _zz_invSub_4 = invSboxRom_166;
      8'b10100111 : _zz_invSub_4 = invSboxRom_167;
      8'b10101000 : _zz_invSub_4 = invSboxRom_168;
      8'b10101001 : _zz_invSub_4 = invSboxRom_169;
      8'b10101010 : _zz_invSub_4 = invSboxRom_170;
      8'b10101011 : _zz_invSub_4 = invSboxRom_171;
      8'b10101100 : _zz_invSub_4 = invSboxRom_172;
      8'b10101101 : _zz_invSub_4 = invSboxRom_173;
      8'b10101110 : _zz_invSub_4 = invSboxRom_174;
      8'b10101111 : _zz_invSub_4 = invSboxRom_175;
      8'b10110000 : _zz_invSub_4 = invSboxRom_176;
      8'b10110001 : _zz_invSub_4 = invSboxRom_177;
      8'b10110010 : _zz_invSub_4 = invSboxRom_178;
      8'b10110011 : _zz_invSub_4 = invSboxRom_179;
      8'b10110100 : _zz_invSub_4 = invSboxRom_180;
      8'b10110101 : _zz_invSub_4 = invSboxRom_181;
      8'b10110110 : _zz_invSub_4 = invSboxRom_182;
      8'b10110111 : _zz_invSub_4 = invSboxRom_183;
      8'b10111000 : _zz_invSub_4 = invSboxRom_184;
      8'b10111001 : _zz_invSub_4 = invSboxRom_185;
      8'b10111010 : _zz_invSub_4 = invSboxRom_186;
      8'b10111011 : _zz_invSub_4 = invSboxRom_187;
      8'b10111100 : _zz_invSub_4 = invSboxRom_188;
      8'b10111101 : _zz_invSub_4 = invSboxRom_189;
      8'b10111110 : _zz_invSub_4 = invSboxRom_190;
      8'b10111111 : _zz_invSub_4 = invSboxRom_191;
      8'b11000000 : _zz_invSub_4 = invSboxRom_192;
      8'b11000001 : _zz_invSub_4 = invSboxRom_193;
      8'b11000010 : _zz_invSub_4 = invSboxRom_194;
      8'b11000011 : _zz_invSub_4 = invSboxRom_195;
      8'b11000100 : _zz_invSub_4 = invSboxRom_196;
      8'b11000101 : _zz_invSub_4 = invSboxRom_197;
      8'b11000110 : _zz_invSub_4 = invSboxRom_198;
      8'b11000111 : _zz_invSub_4 = invSboxRom_199;
      8'b11001000 : _zz_invSub_4 = invSboxRom_200;
      8'b11001001 : _zz_invSub_4 = invSboxRom_201;
      8'b11001010 : _zz_invSub_4 = invSboxRom_202;
      8'b11001011 : _zz_invSub_4 = invSboxRom_203;
      8'b11001100 : _zz_invSub_4 = invSboxRom_204;
      8'b11001101 : _zz_invSub_4 = invSboxRom_205;
      8'b11001110 : _zz_invSub_4 = invSboxRom_206;
      8'b11001111 : _zz_invSub_4 = invSboxRom_207;
      8'b11010000 : _zz_invSub_4 = invSboxRom_208;
      8'b11010001 : _zz_invSub_4 = invSboxRom_209;
      8'b11010010 : _zz_invSub_4 = invSboxRom_210;
      8'b11010011 : _zz_invSub_4 = invSboxRom_211;
      8'b11010100 : _zz_invSub_4 = invSboxRom_212;
      8'b11010101 : _zz_invSub_4 = invSboxRom_213;
      8'b11010110 : _zz_invSub_4 = invSboxRom_214;
      8'b11010111 : _zz_invSub_4 = invSboxRom_215;
      8'b11011000 : _zz_invSub_4 = invSboxRom_216;
      8'b11011001 : _zz_invSub_4 = invSboxRom_217;
      8'b11011010 : _zz_invSub_4 = invSboxRom_218;
      8'b11011011 : _zz_invSub_4 = invSboxRom_219;
      8'b11011100 : _zz_invSub_4 = invSboxRom_220;
      8'b11011101 : _zz_invSub_4 = invSboxRom_221;
      8'b11011110 : _zz_invSub_4 = invSboxRom_222;
      8'b11011111 : _zz_invSub_4 = invSboxRom_223;
      8'b11100000 : _zz_invSub_4 = invSboxRom_224;
      8'b11100001 : _zz_invSub_4 = invSboxRom_225;
      8'b11100010 : _zz_invSub_4 = invSboxRom_226;
      8'b11100011 : _zz_invSub_4 = invSboxRom_227;
      8'b11100100 : _zz_invSub_4 = invSboxRom_228;
      8'b11100101 : _zz_invSub_4 = invSboxRom_229;
      8'b11100110 : _zz_invSub_4 = invSboxRom_230;
      8'b11100111 : _zz_invSub_4 = invSboxRom_231;
      8'b11101000 : _zz_invSub_4 = invSboxRom_232;
      8'b11101001 : _zz_invSub_4 = invSboxRom_233;
      8'b11101010 : _zz_invSub_4 = invSboxRom_234;
      8'b11101011 : _zz_invSub_4 = invSboxRom_235;
      8'b11101100 : _zz_invSub_4 = invSboxRom_236;
      8'b11101101 : _zz_invSub_4 = invSboxRom_237;
      8'b11101110 : _zz_invSub_4 = invSboxRom_238;
      8'b11101111 : _zz_invSub_4 = invSboxRom_239;
      8'b11110000 : _zz_invSub_4 = invSboxRom_240;
      8'b11110001 : _zz_invSub_4 = invSboxRom_241;
      8'b11110010 : _zz_invSub_4 = invSboxRom_242;
      8'b11110011 : _zz_invSub_4 = invSboxRom_243;
      8'b11110100 : _zz_invSub_4 = invSboxRom_244;
      8'b11110101 : _zz_invSub_4 = invSboxRom_245;
      8'b11110110 : _zz_invSub_4 = invSboxRom_246;
      8'b11110111 : _zz_invSub_4 = invSboxRom_247;
      8'b11111000 : _zz_invSub_4 = invSboxRom_248;
      8'b11111001 : _zz_invSub_4 = invSboxRom_249;
      8'b11111010 : _zz_invSub_4 = invSboxRom_250;
      8'b11111011 : _zz_invSub_4 = invSboxRom_251;
      8'b11111100 : _zz_invSub_4 = invSboxRom_252;
      8'b11111101 : _zz_invSub_4 = invSboxRom_253;
      8'b11111110 : _zz_invSub_4 = invSboxRom_254;
      default : _zz_invSub_4 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_5)
      8'b00000000 : _zz_invSub_5 = invSboxRom_0;
      8'b00000001 : _zz_invSub_5 = invSboxRom_1;
      8'b00000010 : _zz_invSub_5 = invSboxRom_2;
      8'b00000011 : _zz_invSub_5 = invSboxRom_3;
      8'b00000100 : _zz_invSub_5 = invSboxRom_4;
      8'b00000101 : _zz_invSub_5 = invSboxRom_5;
      8'b00000110 : _zz_invSub_5 = invSboxRom_6;
      8'b00000111 : _zz_invSub_5 = invSboxRom_7;
      8'b00001000 : _zz_invSub_5 = invSboxRom_8;
      8'b00001001 : _zz_invSub_5 = invSboxRom_9;
      8'b00001010 : _zz_invSub_5 = invSboxRom_10;
      8'b00001011 : _zz_invSub_5 = invSboxRom_11;
      8'b00001100 : _zz_invSub_5 = invSboxRom_12;
      8'b00001101 : _zz_invSub_5 = invSboxRom_13;
      8'b00001110 : _zz_invSub_5 = invSboxRom_14;
      8'b00001111 : _zz_invSub_5 = invSboxRom_15;
      8'b00010000 : _zz_invSub_5 = invSboxRom_16;
      8'b00010001 : _zz_invSub_5 = invSboxRom_17;
      8'b00010010 : _zz_invSub_5 = invSboxRom_18;
      8'b00010011 : _zz_invSub_5 = invSboxRom_19;
      8'b00010100 : _zz_invSub_5 = invSboxRom_20;
      8'b00010101 : _zz_invSub_5 = invSboxRom_21;
      8'b00010110 : _zz_invSub_5 = invSboxRom_22;
      8'b00010111 : _zz_invSub_5 = invSboxRom_23;
      8'b00011000 : _zz_invSub_5 = invSboxRom_24;
      8'b00011001 : _zz_invSub_5 = invSboxRom_25;
      8'b00011010 : _zz_invSub_5 = invSboxRom_26;
      8'b00011011 : _zz_invSub_5 = invSboxRom_27;
      8'b00011100 : _zz_invSub_5 = invSboxRom_28;
      8'b00011101 : _zz_invSub_5 = invSboxRom_29;
      8'b00011110 : _zz_invSub_5 = invSboxRom_30;
      8'b00011111 : _zz_invSub_5 = invSboxRom_31;
      8'b00100000 : _zz_invSub_5 = invSboxRom_32;
      8'b00100001 : _zz_invSub_5 = invSboxRom_33;
      8'b00100010 : _zz_invSub_5 = invSboxRom_34;
      8'b00100011 : _zz_invSub_5 = invSboxRom_35;
      8'b00100100 : _zz_invSub_5 = invSboxRom_36;
      8'b00100101 : _zz_invSub_5 = invSboxRom_37;
      8'b00100110 : _zz_invSub_5 = invSboxRom_38;
      8'b00100111 : _zz_invSub_5 = invSboxRom_39;
      8'b00101000 : _zz_invSub_5 = invSboxRom_40;
      8'b00101001 : _zz_invSub_5 = invSboxRom_41;
      8'b00101010 : _zz_invSub_5 = invSboxRom_42;
      8'b00101011 : _zz_invSub_5 = invSboxRom_43;
      8'b00101100 : _zz_invSub_5 = invSboxRom_44;
      8'b00101101 : _zz_invSub_5 = invSboxRom_45;
      8'b00101110 : _zz_invSub_5 = invSboxRom_46;
      8'b00101111 : _zz_invSub_5 = invSboxRom_47;
      8'b00110000 : _zz_invSub_5 = invSboxRom_48;
      8'b00110001 : _zz_invSub_5 = invSboxRom_49;
      8'b00110010 : _zz_invSub_5 = invSboxRom_50;
      8'b00110011 : _zz_invSub_5 = invSboxRom_51;
      8'b00110100 : _zz_invSub_5 = invSboxRom_52;
      8'b00110101 : _zz_invSub_5 = invSboxRom_53;
      8'b00110110 : _zz_invSub_5 = invSboxRom_54;
      8'b00110111 : _zz_invSub_5 = invSboxRom_55;
      8'b00111000 : _zz_invSub_5 = invSboxRom_56;
      8'b00111001 : _zz_invSub_5 = invSboxRom_57;
      8'b00111010 : _zz_invSub_5 = invSboxRom_58;
      8'b00111011 : _zz_invSub_5 = invSboxRom_59;
      8'b00111100 : _zz_invSub_5 = invSboxRom_60;
      8'b00111101 : _zz_invSub_5 = invSboxRom_61;
      8'b00111110 : _zz_invSub_5 = invSboxRom_62;
      8'b00111111 : _zz_invSub_5 = invSboxRom_63;
      8'b01000000 : _zz_invSub_5 = invSboxRom_64;
      8'b01000001 : _zz_invSub_5 = invSboxRom_65;
      8'b01000010 : _zz_invSub_5 = invSboxRom_66;
      8'b01000011 : _zz_invSub_5 = invSboxRom_67;
      8'b01000100 : _zz_invSub_5 = invSboxRom_68;
      8'b01000101 : _zz_invSub_5 = invSboxRom_69;
      8'b01000110 : _zz_invSub_5 = invSboxRom_70;
      8'b01000111 : _zz_invSub_5 = invSboxRom_71;
      8'b01001000 : _zz_invSub_5 = invSboxRom_72;
      8'b01001001 : _zz_invSub_5 = invSboxRom_73;
      8'b01001010 : _zz_invSub_5 = invSboxRom_74;
      8'b01001011 : _zz_invSub_5 = invSboxRom_75;
      8'b01001100 : _zz_invSub_5 = invSboxRom_76;
      8'b01001101 : _zz_invSub_5 = invSboxRom_77;
      8'b01001110 : _zz_invSub_5 = invSboxRom_78;
      8'b01001111 : _zz_invSub_5 = invSboxRom_79;
      8'b01010000 : _zz_invSub_5 = invSboxRom_80;
      8'b01010001 : _zz_invSub_5 = invSboxRom_81;
      8'b01010010 : _zz_invSub_5 = invSboxRom_82;
      8'b01010011 : _zz_invSub_5 = invSboxRom_83;
      8'b01010100 : _zz_invSub_5 = invSboxRom_84;
      8'b01010101 : _zz_invSub_5 = invSboxRom_85;
      8'b01010110 : _zz_invSub_5 = invSboxRom_86;
      8'b01010111 : _zz_invSub_5 = invSboxRom_87;
      8'b01011000 : _zz_invSub_5 = invSboxRom_88;
      8'b01011001 : _zz_invSub_5 = invSboxRom_89;
      8'b01011010 : _zz_invSub_5 = invSboxRom_90;
      8'b01011011 : _zz_invSub_5 = invSboxRom_91;
      8'b01011100 : _zz_invSub_5 = invSboxRom_92;
      8'b01011101 : _zz_invSub_5 = invSboxRom_93;
      8'b01011110 : _zz_invSub_5 = invSboxRom_94;
      8'b01011111 : _zz_invSub_5 = invSboxRom_95;
      8'b01100000 : _zz_invSub_5 = invSboxRom_96;
      8'b01100001 : _zz_invSub_5 = invSboxRom_97;
      8'b01100010 : _zz_invSub_5 = invSboxRom_98;
      8'b01100011 : _zz_invSub_5 = invSboxRom_99;
      8'b01100100 : _zz_invSub_5 = invSboxRom_100;
      8'b01100101 : _zz_invSub_5 = invSboxRom_101;
      8'b01100110 : _zz_invSub_5 = invSboxRom_102;
      8'b01100111 : _zz_invSub_5 = invSboxRom_103;
      8'b01101000 : _zz_invSub_5 = invSboxRom_104;
      8'b01101001 : _zz_invSub_5 = invSboxRom_105;
      8'b01101010 : _zz_invSub_5 = invSboxRom_106;
      8'b01101011 : _zz_invSub_5 = invSboxRom_107;
      8'b01101100 : _zz_invSub_5 = invSboxRom_108;
      8'b01101101 : _zz_invSub_5 = invSboxRom_109;
      8'b01101110 : _zz_invSub_5 = invSboxRom_110;
      8'b01101111 : _zz_invSub_5 = invSboxRom_111;
      8'b01110000 : _zz_invSub_5 = invSboxRom_112;
      8'b01110001 : _zz_invSub_5 = invSboxRom_113;
      8'b01110010 : _zz_invSub_5 = invSboxRom_114;
      8'b01110011 : _zz_invSub_5 = invSboxRom_115;
      8'b01110100 : _zz_invSub_5 = invSboxRom_116;
      8'b01110101 : _zz_invSub_5 = invSboxRom_117;
      8'b01110110 : _zz_invSub_5 = invSboxRom_118;
      8'b01110111 : _zz_invSub_5 = invSboxRom_119;
      8'b01111000 : _zz_invSub_5 = invSboxRom_120;
      8'b01111001 : _zz_invSub_5 = invSboxRom_121;
      8'b01111010 : _zz_invSub_5 = invSboxRom_122;
      8'b01111011 : _zz_invSub_5 = invSboxRom_123;
      8'b01111100 : _zz_invSub_5 = invSboxRom_124;
      8'b01111101 : _zz_invSub_5 = invSboxRom_125;
      8'b01111110 : _zz_invSub_5 = invSboxRom_126;
      8'b01111111 : _zz_invSub_5 = invSboxRom_127;
      8'b10000000 : _zz_invSub_5 = invSboxRom_128;
      8'b10000001 : _zz_invSub_5 = invSboxRom_129;
      8'b10000010 : _zz_invSub_5 = invSboxRom_130;
      8'b10000011 : _zz_invSub_5 = invSboxRom_131;
      8'b10000100 : _zz_invSub_5 = invSboxRom_132;
      8'b10000101 : _zz_invSub_5 = invSboxRom_133;
      8'b10000110 : _zz_invSub_5 = invSboxRom_134;
      8'b10000111 : _zz_invSub_5 = invSboxRom_135;
      8'b10001000 : _zz_invSub_5 = invSboxRom_136;
      8'b10001001 : _zz_invSub_5 = invSboxRom_137;
      8'b10001010 : _zz_invSub_5 = invSboxRom_138;
      8'b10001011 : _zz_invSub_5 = invSboxRom_139;
      8'b10001100 : _zz_invSub_5 = invSboxRom_140;
      8'b10001101 : _zz_invSub_5 = invSboxRom_141;
      8'b10001110 : _zz_invSub_5 = invSboxRom_142;
      8'b10001111 : _zz_invSub_5 = invSboxRom_143;
      8'b10010000 : _zz_invSub_5 = invSboxRom_144;
      8'b10010001 : _zz_invSub_5 = invSboxRom_145;
      8'b10010010 : _zz_invSub_5 = invSboxRom_146;
      8'b10010011 : _zz_invSub_5 = invSboxRom_147;
      8'b10010100 : _zz_invSub_5 = invSboxRom_148;
      8'b10010101 : _zz_invSub_5 = invSboxRom_149;
      8'b10010110 : _zz_invSub_5 = invSboxRom_150;
      8'b10010111 : _zz_invSub_5 = invSboxRom_151;
      8'b10011000 : _zz_invSub_5 = invSboxRom_152;
      8'b10011001 : _zz_invSub_5 = invSboxRom_153;
      8'b10011010 : _zz_invSub_5 = invSboxRom_154;
      8'b10011011 : _zz_invSub_5 = invSboxRom_155;
      8'b10011100 : _zz_invSub_5 = invSboxRom_156;
      8'b10011101 : _zz_invSub_5 = invSboxRom_157;
      8'b10011110 : _zz_invSub_5 = invSboxRom_158;
      8'b10011111 : _zz_invSub_5 = invSboxRom_159;
      8'b10100000 : _zz_invSub_5 = invSboxRom_160;
      8'b10100001 : _zz_invSub_5 = invSboxRom_161;
      8'b10100010 : _zz_invSub_5 = invSboxRom_162;
      8'b10100011 : _zz_invSub_5 = invSboxRom_163;
      8'b10100100 : _zz_invSub_5 = invSboxRom_164;
      8'b10100101 : _zz_invSub_5 = invSboxRom_165;
      8'b10100110 : _zz_invSub_5 = invSboxRom_166;
      8'b10100111 : _zz_invSub_5 = invSboxRom_167;
      8'b10101000 : _zz_invSub_5 = invSboxRom_168;
      8'b10101001 : _zz_invSub_5 = invSboxRom_169;
      8'b10101010 : _zz_invSub_5 = invSboxRom_170;
      8'b10101011 : _zz_invSub_5 = invSboxRom_171;
      8'b10101100 : _zz_invSub_5 = invSboxRom_172;
      8'b10101101 : _zz_invSub_5 = invSboxRom_173;
      8'b10101110 : _zz_invSub_5 = invSboxRom_174;
      8'b10101111 : _zz_invSub_5 = invSboxRom_175;
      8'b10110000 : _zz_invSub_5 = invSboxRom_176;
      8'b10110001 : _zz_invSub_5 = invSboxRom_177;
      8'b10110010 : _zz_invSub_5 = invSboxRom_178;
      8'b10110011 : _zz_invSub_5 = invSboxRom_179;
      8'b10110100 : _zz_invSub_5 = invSboxRom_180;
      8'b10110101 : _zz_invSub_5 = invSboxRom_181;
      8'b10110110 : _zz_invSub_5 = invSboxRom_182;
      8'b10110111 : _zz_invSub_5 = invSboxRom_183;
      8'b10111000 : _zz_invSub_5 = invSboxRom_184;
      8'b10111001 : _zz_invSub_5 = invSboxRom_185;
      8'b10111010 : _zz_invSub_5 = invSboxRom_186;
      8'b10111011 : _zz_invSub_5 = invSboxRom_187;
      8'b10111100 : _zz_invSub_5 = invSboxRom_188;
      8'b10111101 : _zz_invSub_5 = invSboxRom_189;
      8'b10111110 : _zz_invSub_5 = invSboxRom_190;
      8'b10111111 : _zz_invSub_5 = invSboxRom_191;
      8'b11000000 : _zz_invSub_5 = invSboxRom_192;
      8'b11000001 : _zz_invSub_5 = invSboxRom_193;
      8'b11000010 : _zz_invSub_5 = invSboxRom_194;
      8'b11000011 : _zz_invSub_5 = invSboxRom_195;
      8'b11000100 : _zz_invSub_5 = invSboxRom_196;
      8'b11000101 : _zz_invSub_5 = invSboxRom_197;
      8'b11000110 : _zz_invSub_5 = invSboxRom_198;
      8'b11000111 : _zz_invSub_5 = invSboxRom_199;
      8'b11001000 : _zz_invSub_5 = invSboxRom_200;
      8'b11001001 : _zz_invSub_5 = invSboxRom_201;
      8'b11001010 : _zz_invSub_5 = invSboxRom_202;
      8'b11001011 : _zz_invSub_5 = invSboxRom_203;
      8'b11001100 : _zz_invSub_5 = invSboxRom_204;
      8'b11001101 : _zz_invSub_5 = invSboxRom_205;
      8'b11001110 : _zz_invSub_5 = invSboxRom_206;
      8'b11001111 : _zz_invSub_5 = invSboxRom_207;
      8'b11010000 : _zz_invSub_5 = invSboxRom_208;
      8'b11010001 : _zz_invSub_5 = invSboxRom_209;
      8'b11010010 : _zz_invSub_5 = invSboxRom_210;
      8'b11010011 : _zz_invSub_5 = invSboxRom_211;
      8'b11010100 : _zz_invSub_5 = invSboxRom_212;
      8'b11010101 : _zz_invSub_5 = invSboxRom_213;
      8'b11010110 : _zz_invSub_5 = invSboxRom_214;
      8'b11010111 : _zz_invSub_5 = invSboxRom_215;
      8'b11011000 : _zz_invSub_5 = invSboxRom_216;
      8'b11011001 : _zz_invSub_5 = invSboxRom_217;
      8'b11011010 : _zz_invSub_5 = invSboxRom_218;
      8'b11011011 : _zz_invSub_5 = invSboxRom_219;
      8'b11011100 : _zz_invSub_5 = invSboxRom_220;
      8'b11011101 : _zz_invSub_5 = invSboxRom_221;
      8'b11011110 : _zz_invSub_5 = invSboxRom_222;
      8'b11011111 : _zz_invSub_5 = invSboxRom_223;
      8'b11100000 : _zz_invSub_5 = invSboxRom_224;
      8'b11100001 : _zz_invSub_5 = invSboxRom_225;
      8'b11100010 : _zz_invSub_5 = invSboxRom_226;
      8'b11100011 : _zz_invSub_5 = invSboxRom_227;
      8'b11100100 : _zz_invSub_5 = invSboxRom_228;
      8'b11100101 : _zz_invSub_5 = invSboxRom_229;
      8'b11100110 : _zz_invSub_5 = invSboxRom_230;
      8'b11100111 : _zz_invSub_5 = invSboxRom_231;
      8'b11101000 : _zz_invSub_5 = invSboxRom_232;
      8'b11101001 : _zz_invSub_5 = invSboxRom_233;
      8'b11101010 : _zz_invSub_5 = invSboxRom_234;
      8'b11101011 : _zz_invSub_5 = invSboxRom_235;
      8'b11101100 : _zz_invSub_5 = invSboxRom_236;
      8'b11101101 : _zz_invSub_5 = invSboxRom_237;
      8'b11101110 : _zz_invSub_5 = invSboxRom_238;
      8'b11101111 : _zz_invSub_5 = invSboxRom_239;
      8'b11110000 : _zz_invSub_5 = invSboxRom_240;
      8'b11110001 : _zz_invSub_5 = invSboxRom_241;
      8'b11110010 : _zz_invSub_5 = invSboxRom_242;
      8'b11110011 : _zz_invSub_5 = invSboxRom_243;
      8'b11110100 : _zz_invSub_5 = invSboxRom_244;
      8'b11110101 : _zz_invSub_5 = invSboxRom_245;
      8'b11110110 : _zz_invSub_5 = invSboxRom_246;
      8'b11110111 : _zz_invSub_5 = invSboxRom_247;
      8'b11111000 : _zz_invSub_5 = invSboxRom_248;
      8'b11111001 : _zz_invSub_5 = invSboxRom_249;
      8'b11111010 : _zz_invSub_5 = invSboxRom_250;
      8'b11111011 : _zz_invSub_5 = invSboxRom_251;
      8'b11111100 : _zz_invSub_5 = invSboxRom_252;
      8'b11111101 : _zz_invSub_5 = invSboxRom_253;
      8'b11111110 : _zz_invSub_5 = invSboxRom_254;
      default : _zz_invSub_5 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_6)
      8'b00000000 : _zz_invSub_6 = invSboxRom_0;
      8'b00000001 : _zz_invSub_6 = invSboxRom_1;
      8'b00000010 : _zz_invSub_6 = invSboxRom_2;
      8'b00000011 : _zz_invSub_6 = invSboxRom_3;
      8'b00000100 : _zz_invSub_6 = invSboxRom_4;
      8'b00000101 : _zz_invSub_6 = invSboxRom_5;
      8'b00000110 : _zz_invSub_6 = invSboxRom_6;
      8'b00000111 : _zz_invSub_6 = invSboxRom_7;
      8'b00001000 : _zz_invSub_6 = invSboxRom_8;
      8'b00001001 : _zz_invSub_6 = invSboxRom_9;
      8'b00001010 : _zz_invSub_6 = invSboxRom_10;
      8'b00001011 : _zz_invSub_6 = invSboxRom_11;
      8'b00001100 : _zz_invSub_6 = invSboxRom_12;
      8'b00001101 : _zz_invSub_6 = invSboxRom_13;
      8'b00001110 : _zz_invSub_6 = invSboxRom_14;
      8'b00001111 : _zz_invSub_6 = invSboxRom_15;
      8'b00010000 : _zz_invSub_6 = invSboxRom_16;
      8'b00010001 : _zz_invSub_6 = invSboxRom_17;
      8'b00010010 : _zz_invSub_6 = invSboxRom_18;
      8'b00010011 : _zz_invSub_6 = invSboxRom_19;
      8'b00010100 : _zz_invSub_6 = invSboxRom_20;
      8'b00010101 : _zz_invSub_6 = invSboxRom_21;
      8'b00010110 : _zz_invSub_6 = invSboxRom_22;
      8'b00010111 : _zz_invSub_6 = invSboxRom_23;
      8'b00011000 : _zz_invSub_6 = invSboxRom_24;
      8'b00011001 : _zz_invSub_6 = invSboxRom_25;
      8'b00011010 : _zz_invSub_6 = invSboxRom_26;
      8'b00011011 : _zz_invSub_6 = invSboxRom_27;
      8'b00011100 : _zz_invSub_6 = invSboxRom_28;
      8'b00011101 : _zz_invSub_6 = invSboxRom_29;
      8'b00011110 : _zz_invSub_6 = invSboxRom_30;
      8'b00011111 : _zz_invSub_6 = invSboxRom_31;
      8'b00100000 : _zz_invSub_6 = invSboxRom_32;
      8'b00100001 : _zz_invSub_6 = invSboxRom_33;
      8'b00100010 : _zz_invSub_6 = invSboxRom_34;
      8'b00100011 : _zz_invSub_6 = invSboxRom_35;
      8'b00100100 : _zz_invSub_6 = invSboxRom_36;
      8'b00100101 : _zz_invSub_6 = invSboxRom_37;
      8'b00100110 : _zz_invSub_6 = invSboxRom_38;
      8'b00100111 : _zz_invSub_6 = invSboxRom_39;
      8'b00101000 : _zz_invSub_6 = invSboxRom_40;
      8'b00101001 : _zz_invSub_6 = invSboxRom_41;
      8'b00101010 : _zz_invSub_6 = invSboxRom_42;
      8'b00101011 : _zz_invSub_6 = invSboxRom_43;
      8'b00101100 : _zz_invSub_6 = invSboxRom_44;
      8'b00101101 : _zz_invSub_6 = invSboxRom_45;
      8'b00101110 : _zz_invSub_6 = invSboxRom_46;
      8'b00101111 : _zz_invSub_6 = invSboxRom_47;
      8'b00110000 : _zz_invSub_6 = invSboxRom_48;
      8'b00110001 : _zz_invSub_6 = invSboxRom_49;
      8'b00110010 : _zz_invSub_6 = invSboxRom_50;
      8'b00110011 : _zz_invSub_6 = invSboxRom_51;
      8'b00110100 : _zz_invSub_6 = invSboxRom_52;
      8'b00110101 : _zz_invSub_6 = invSboxRom_53;
      8'b00110110 : _zz_invSub_6 = invSboxRom_54;
      8'b00110111 : _zz_invSub_6 = invSboxRom_55;
      8'b00111000 : _zz_invSub_6 = invSboxRom_56;
      8'b00111001 : _zz_invSub_6 = invSboxRom_57;
      8'b00111010 : _zz_invSub_6 = invSboxRom_58;
      8'b00111011 : _zz_invSub_6 = invSboxRom_59;
      8'b00111100 : _zz_invSub_6 = invSboxRom_60;
      8'b00111101 : _zz_invSub_6 = invSboxRom_61;
      8'b00111110 : _zz_invSub_6 = invSboxRom_62;
      8'b00111111 : _zz_invSub_6 = invSboxRom_63;
      8'b01000000 : _zz_invSub_6 = invSboxRom_64;
      8'b01000001 : _zz_invSub_6 = invSboxRom_65;
      8'b01000010 : _zz_invSub_6 = invSboxRom_66;
      8'b01000011 : _zz_invSub_6 = invSboxRom_67;
      8'b01000100 : _zz_invSub_6 = invSboxRom_68;
      8'b01000101 : _zz_invSub_6 = invSboxRom_69;
      8'b01000110 : _zz_invSub_6 = invSboxRom_70;
      8'b01000111 : _zz_invSub_6 = invSboxRom_71;
      8'b01001000 : _zz_invSub_6 = invSboxRom_72;
      8'b01001001 : _zz_invSub_6 = invSboxRom_73;
      8'b01001010 : _zz_invSub_6 = invSboxRom_74;
      8'b01001011 : _zz_invSub_6 = invSboxRom_75;
      8'b01001100 : _zz_invSub_6 = invSboxRom_76;
      8'b01001101 : _zz_invSub_6 = invSboxRom_77;
      8'b01001110 : _zz_invSub_6 = invSboxRom_78;
      8'b01001111 : _zz_invSub_6 = invSboxRom_79;
      8'b01010000 : _zz_invSub_6 = invSboxRom_80;
      8'b01010001 : _zz_invSub_6 = invSboxRom_81;
      8'b01010010 : _zz_invSub_6 = invSboxRom_82;
      8'b01010011 : _zz_invSub_6 = invSboxRom_83;
      8'b01010100 : _zz_invSub_6 = invSboxRom_84;
      8'b01010101 : _zz_invSub_6 = invSboxRom_85;
      8'b01010110 : _zz_invSub_6 = invSboxRom_86;
      8'b01010111 : _zz_invSub_6 = invSboxRom_87;
      8'b01011000 : _zz_invSub_6 = invSboxRom_88;
      8'b01011001 : _zz_invSub_6 = invSboxRom_89;
      8'b01011010 : _zz_invSub_6 = invSboxRom_90;
      8'b01011011 : _zz_invSub_6 = invSboxRom_91;
      8'b01011100 : _zz_invSub_6 = invSboxRom_92;
      8'b01011101 : _zz_invSub_6 = invSboxRom_93;
      8'b01011110 : _zz_invSub_6 = invSboxRom_94;
      8'b01011111 : _zz_invSub_6 = invSboxRom_95;
      8'b01100000 : _zz_invSub_6 = invSboxRom_96;
      8'b01100001 : _zz_invSub_6 = invSboxRom_97;
      8'b01100010 : _zz_invSub_6 = invSboxRom_98;
      8'b01100011 : _zz_invSub_6 = invSboxRom_99;
      8'b01100100 : _zz_invSub_6 = invSboxRom_100;
      8'b01100101 : _zz_invSub_6 = invSboxRom_101;
      8'b01100110 : _zz_invSub_6 = invSboxRom_102;
      8'b01100111 : _zz_invSub_6 = invSboxRom_103;
      8'b01101000 : _zz_invSub_6 = invSboxRom_104;
      8'b01101001 : _zz_invSub_6 = invSboxRom_105;
      8'b01101010 : _zz_invSub_6 = invSboxRom_106;
      8'b01101011 : _zz_invSub_6 = invSboxRom_107;
      8'b01101100 : _zz_invSub_6 = invSboxRom_108;
      8'b01101101 : _zz_invSub_6 = invSboxRom_109;
      8'b01101110 : _zz_invSub_6 = invSboxRom_110;
      8'b01101111 : _zz_invSub_6 = invSboxRom_111;
      8'b01110000 : _zz_invSub_6 = invSboxRom_112;
      8'b01110001 : _zz_invSub_6 = invSboxRom_113;
      8'b01110010 : _zz_invSub_6 = invSboxRom_114;
      8'b01110011 : _zz_invSub_6 = invSboxRom_115;
      8'b01110100 : _zz_invSub_6 = invSboxRom_116;
      8'b01110101 : _zz_invSub_6 = invSboxRom_117;
      8'b01110110 : _zz_invSub_6 = invSboxRom_118;
      8'b01110111 : _zz_invSub_6 = invSboxRom_119;
      8'b01111000 : _zz_invSub_6 = invSboxRom_120;
      8'b01111001 : _zz_invSub_6 = invSboxRom_121;
      8'b01111010 : _zz_invSub_6 = invSboxRom_122;
      8'b01111011 : _zz_invSub_6 = invSboxRom_123;
      8'b01111100 : _zz_invSub_6 = invSboxRom_124;
      8'b01111101 : _zz_invSub_6 = invSboxRom_125;
      8'b01111110 : _zz_invSub_6 = invSboxRom_126;
      8'b01111111 : _zz_invSub_6 = invSboxRom_127;
      8'b10000000 : _zz_invSub_6 = invSboxRom_128;
      8'b10000001 : _zz_invSub_6 = invSboxRom_129;
      8'b10000010 : _zz_invSub_6 = invSboxRom_130;
      8'b10000011 : _zz_invSub_6 = invSboxRom_131;
      8'b10000100 : _zz_invSub_6 = invSboxRom_132;
      8'b10000101 : _zz_invSub_6 = invSboxRom_133;
      8'b10000110 : _zz_invSub_6 = invSboxRom_134;
      8'b10000111 : _zz_invSub_6 = invSboxRom_135;
      8'b10001000 : _zz_invSub_6 = invSboxRom_136;
      8'b10001001 : _zz_invSub_6 = invSboxRom_137;
      8'b10001010 : _zz_invSub_6 = invSboxRom_138;
      8'b10001011 : _zz_invSub_6 = invSboxRom_139;
      8'b10001100 : _zz_invSub_6 = invSboxRom_140;
      8'b10001101 : _zz_invSub_6 = invSboxRom_141;
      8'b10001110 : _zz_invSub_6 = invSboxRom_142;
      8'b10001111 : _zz_invSub_6 = invSboxRom_143;
      8'b10010000 : _zz_invSub_6 = invSboxRom_144;
      8'b10010001 : _zz_invSub_6 = invSboxRom_145;
      8'b10010010 : _zz_invSub_6 = invSboxRom_146;
      8'b10010011 : _zz_invSub_6 = invSboxRom_147;
      8'b10010100 : _zz_invSub_6 = invSboxRom_148;
      8'b10010101 : _zz_invSub_6 = invSboxRom_149;
      8'b10010110 : _zz_invSub_6 = invSboxRom_150;
      8'b10010111 : _zz_invSub_6 = invSboxRom_151;
      8'b10011000 : _zz_invSub_6 = invSboxRom_152;
      8'b10011001 : _zz_invSub_6 = invSboxRom_153;
      8'b10011010 : _zz_invSub_6 = invSboxRom_154;
      8'b10011011 : _zz_invSub_6 = invSboxRom_155;
      8'b10011100 : _zz_invSub_6 = invSboxRom_156;
      8'b10011101 : _zz_invSub_6 = invSboxRom_157;
      8'b10011110 : _zz_invSub_6 = invSboxRom_158;
      8'b10011111 : _zz_invSub_6 = invSboxRom_159;
      8'b10100000 : _zz_invSub_6 = invSboxRom_160;
      8'b10100001 : _zz_invSub_6 = invSboxRom_161;
      8'b10100010 : _zz_invSub_6 = invSboxRom_162;
      8'b10100011 : _zz_invSub_6 = invSboxRom_163;
      8'b10100100 : _zz_invSub_6 = invSboxRom_164;
      8'b10100101 : _zz_invSub_6 = invSboxRom_165;
      8'b10100110 : _zz_invSub_6 = invSboxRom_166;
      8'b10100111 : _zz_invSub_6 = invSboxRom_167;
      8'b10101000 : _zz_invSub_6 = invSboxRom_168;
      8'b10101001 : _zz_invSub_6 = invSboxRom_169;
      8'b10101010 : _zz_invSub_6 = invSboxRom_170;
      8'b10101011 : _zz_invSub_6 = invSboxRom_171;
      8'b10101100 : _zz_invSub_6 = invSboxRom_172;
      8'b10101101 : _zz_invSub_6 = invSboxRom_173;
      8'b10101110 : _zz_invSub_6 = invSboxRom_174;
      8'b10101111 : _zz_invSub_6 = invSboxRom_175;
      8'b10110000 : _zz_invSub_6 = invSboxRom_176;
      8'b10110001 : _zz_invSub_6 = invSboxRom_177;
      8'b10110010 : _zz_invSub_6 = invSboxRom_178;
      8'b10110011 : _zz_invSub_6 = invSboxRom_179;
      8'b10110100 : _zz_invSub_6 = invSboxRom_180;
      8'b10110101 : _zz_invSub_6 = invSboxRom_181;
      8'b10110110 : _zz_invSub_6 = invSboxRom_182;
      8'b10110111 : _zz_invSub_6 = invSboxRom_183;
      8'b10111000 : _zz_invSub_6 = invSboxRom_184;
      8'b10111001 : _zz_invSub_6 = invSboxRom_185;
      8'b10111010 : _zz_invSub_6 = invSboxRom_186;
      8'b10111011 : _zz_invSub_6 = invSboxRom_187;
      8'b10111100 : _zz_invSub_6 = invSboxRom_188;
      8'b10111101 : _zz_invSub_6 = invSboxRom_189;
      8'b10111110 : _zz_invSub_6 = invSboxRom_190;
      8'b10111111 : _zz_invSub_6 = invSboxRom_191;
      8'b11000000 : _zz_invSub_6 = invSboxRom_192;
      8'b11000001 : _zz_invSub_6 = invSboxRom_193;
      8'b11000010 : _zz_invSub_6 = invSboxRom_194;
      8'b11000011 : _zz_invSub_6 = invSboxRom_195;
      8'b11000100 : _zz_invSub_6 = invSboxRom_196;
      8'b11000101 : _zz_invSub_6 = invSboxRom_197;
      8'b11000110 : _zz_invSub_6 = invSboxRom_198;
      8'b11000111 : _zz_invSub_6 = invSboxRom_199;
      8'b11001000 : _zz_invSub_6 = invSboxRom_200;
      8'b11001001 : _zz_invSub_6 = invSboxRom_201;
      8'b11001010 : _zz_invSub_6 = invSboxRom_202;
      8'b11001011 : _zz_invSub_6 = invSboxRom_203;
      8'b11001100 : _zz_invSub_6 = invSboxRom_204;
      8'b11001101 : _zz_invSub_6 = invSboxRom_205;
      8'b11001110 : _zz_invSub_6 = invSboxRom_206;
      8'b11001111 : _zz_invSub_6 = invSboxRom_207;
      8'b11010000 : _zz_invSub_6 = invSboxRom_208;
      8'b11010001 : _zz_invSub_6 = invSboxRom_209;
      8'b11010010 : _zz_invSub_6 = invSboxRom_210;
      8'b11010011 : _zz_invSub_6 = invSboxRom_211;
      8'b11010100 : _zz_invSub_6 = invSboxRom_212;
      8'b11010101 : _zz_invSub_6 = invSboxRom_213;
      8'b11010110 : _zz_invSub_6 = invSboxRom_214;
      8'b11010111 : _zz_invSub_6 = invSboxRom_215;
      8'b11011000 : _zz_invSub_6 = invSboxRom_216;
      8'b11011001 : _zz_invSub_6 = invSboxRom_217;
      8'b11011010 : _zz_invSub_6 = invSboxRom_218;
      8'b11011011 : _zz_invSub_6 = invSboxRom_219;
      8'b11011100 : _zz_invSub_6 = invSboxRom_220;
      8'b11011101 : _zz_invSub_6 = invSboxRom_221;
      8'b11011110 : _zz_invSub_6 = invSboxRom_222;
      8'b11011111 : _zz_invSub_6 = invSboxRom_223;
      8'b11100000 : _zz_invSub_6 = invSboxRom_224;
      8'b11100001 : _zz_invSub_6 = invSboxRom_225;
      8'b11100010 : _zz_invSub_6 = invSboxRom_226;
      8'b11100011 : _zz_invSub_6 = invSboxRom_227;
      8'b11100100 : _zz_invSub_6 = invSboxRom_228;
      8'b11100101 : _zz_invSub_6 = invSboxRom_229;
      8'b11100110 : _zz_invSub_6 = invSboxRom_230;
      8'b11100111 : _zz_invSub_6 = invSboxRom_231;
      8'b11101000 : _zz_invSub_6 = invSboxRom_232;
      8'b11101001 : _zz_invSub_6 = invSboxRom_233;
      8'b11101010 : _zz_invSub_6 = invSboxRom_234;
      8'b11101011 : _zz_invSub_6 = invSboxRom_235;
      8'b11101100 : _zz_invSub_6 = invSboxRom_236;
      8'b11101101 : _zz_invSub_6 = invSboxRom_237;
      8'b11101110 : _zz_invSub_6 = invSboxRom_238;
      8'b11101111 : _zz_invSub_6 = invSboxRom_239;
      8'b11110000 : _zz_invSub_6 = invSboxRom_240;
      8'b11110001 : _zz_invSub_6 = invSboxRom_241;
      8'b11110010 : _zz_invSub_6 = invSboxRom_242;
      8'b11110011 : _zz_invSub_6 = invSboxRom_243;
      8'b11110100 : _zz_invSub_6 = invSboxRom_244;
      8'b11110101 : _zz_invSub_6 = invSboxRom_245;
      8'b11110110 : _zz_invSub_6 = invSboxRom_246;
      8'b11110111 : _zz_invSub_6 = invSboxRom_247;
      8'b11111000 : _zz_invSub_6 = invSboxRom_248;
      8'b11111001 : _zz_invSub_6 = invSboxRom_249;
      8'b11111010 : _zz_invSub_6 = invSboxRom_250;
      8'b11111011 : _zz_invSub_6 = invSboxRom_251;
      8'b11111100 : _zz_invSub_6 = invSboxRom_252;
      8'b11111101 : _zz_invSub_6 = invSboxRom_253;
      8'b11111110 : _zz_invSub_6 = invSboxRom_254;
      default : _zz_invSub_6 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_7)
      8'b00000000 : _zz_invSub_7 = invSboxRom_0;
      8'b00000001 : _zz_invSub_7 = invSboxRom_1;
      8'b00000010 : _zz_invSub_7 = invSboxRom_2;
      8'b00000011 : _zz_invSub_7 = invSboxRom_3;
      8'b00000100 : _zz_invSub_7 = invSboxRom_4;
      8'b00000101 : _zz_invSub_7 = invSboxRom_5;
      8'b00000110 : _zz_invSub_7 = invSboxRom_6;
      8'b00000111 : _zz_invSub_7 = invSboxRom_7;
      8'b00001000 : _zz_invSub_7 = invSboxRom_8;
      8'b00001001 : _zz_invSub_7 = invSboxRom_9;
      8'b00001010 : _zz_invSub_7 = invSboxRom_10;
      8'b00001011 : _zz_invSub_7 = invSboxRom_11;
      8'b00001100 : _zz_invSub_7 = invSboxRom_12;
      8'b00001101 : _zz_invSub_7 = invSboxRom_13;
      8'b00001110 : _zz_invSub_7 = invSboxRom_14;
      8'b00001111 : _zz_invSub_7 = invSboxRom_15;
      8'b00010000 : _zz_invSub_7 = invSboxRom_16;
      8'b00010001 : _zz_invSub_7 = invSboxRom_17;
      8'b00010010 : _zz_invSub_7 = invSboxRom_18;
      8'b00010011 : _zz_invSub_7 = invSboxRom_19;
      8'b00010100 : _zz_invSub_7 = invSboxRom_20;
      8'b00010101 : _zz_invSub_7 = invSboxRom_21;
      8'b00010110 : _zz_invSub_7 = invSboxRom_22;
      8'b00010111 : _zz_invSub_7 = invSboxRom_23;
      8'b00011000 : _zz_invSub_7 = invSboxRom_24;
      8'b00011001 : _zz_invSub_7 = invSboxRom_25;
      8'b00011010 : _zz_invSub_7 = invSboxRom_26;
      8'b00011011 : _zz_invSub_7 = invSboxRom_27;
      8'b00011100 : _zz_invSub_7 = invSboxRom_28;
      8'b00011101 : _zz_invSub_7 = invSboxRom_29;
      8'b00011110 : _zz_invSub_7 = invSboxRom_30;
      8'b00011111 : _zz_invSub_7 = invSboxRom_31;
      8'b00100000 : _zz_invSub_7 = invSboxRom_32;
      8'b00100001 : _zz_invSub_7 = invSboxRom_33;
      8'b00100010 : _zz_invSub_7 = invSboxRom_34;
      8'b00100011 : _zz_invSub_7 = invSboxRom_35;
      8'b00100100 : _zz_invSub_7 = invSboxRom_36;
      8'b00100101 : _zz_invSub_7 = invSboxRom_37;
      8'b00100110 : _zz_invSub_7 = invSboxRom_38;
      8'b00100111 : _zz_invSub_7 = invSboxRom_39;
      8'b00101000 : _zz_invSub_7 = invSboxRom_40;
      8'b00101001 : _zz_invSub_7 = invSboxRom_41;
      8'b00101010 : _zz_invSub_7 = invSboxRom_42;
      8'b00101011 : _zz_invSub_7 = invSboxRom_43;
      8'b00101100 : _zz_invSub_7 = invSboxRom_44;
      8'b00101101 : _zz_invSub_7 = invSboxRom_45;
      8'b00101110 : _zz_invSub_7 = invSboxRom_46;
      8'b00101111 : _zz_invSub_7 = invSboxRom_47;
      8'b00110000 : _zz_invSub_7 = invSboxRom_48;
      8'b00110001 : _zz_invSub_7 = invSboxRom_49;
      8'b00110010 : _zz_invSub_7 = invSboxRom_50;
      8'b00110011 : _zz_invSub_7 = invSboxRom_51;
      8'b00110100 : _zz_invSub_7 = invSboxRom_52;
      8'b00110101 : _zz_invSub_7 = invSboxRom_53;
      8'b00110110 : _zz_invSub_7 = invSboxRom_54;
      8'b00110111 : _zz_invSub_7 = invSboxRom_55;
      8'b00111000 : _zz_invSub_7 = invSboxRom_56;
      8'b00111001 : _zz_invSub_7 = invSboxRom_57;
      8'b00111010 : _zz_invSub_7 = invSboxRom_58;
      8'b00111011 : _zz_invSub_7 = invSboxRom_59;
      8'b00111100 : _zz_invSub_7 = invSboxRom_60;
      8'b00111101 : _zz_invSub_7 = invSboxRom_61;
      8'b00111110 : _zz_invSub_7 = invSboxRom_62;
      8'b00111111 : _zz_invSub_7 = invSboxRom_63;
      8'b01000000 : _zz_invSub_7 = invSboxRom_64;
      8'b01000001 : _zz_invSub_7 = invSboxRom_65;
      8'b01000010 : _zz_invSub_7 = invSboxRom_66;
      8'b01000011 : _zz_invSub_7 = invSboxRom_67;
      8'b01000100 : _zz_invSub_7 = invSboxRom_68;
      8'b01000101 : _zz_invSub_7 = invSboxRom_69;
      8'b01000110 : _zz_invSub_7 = invSboxRom_70;
      8'b01000111 : _zz_invSub_7 = invSboxRom_71;
      8'b01001000 : _zz_invSub_7 = invSboxRom_72;
      8'b01001001 : _zz_invSub_7 = invSboxRom_73;
      8'b01001010 : _zz_invSub_7 = invSboxRom_74;
      8'b01001011 : _zz_invSub_7 = invSboxRom_75;
      8'b01001100 : _zz_invSub_7 = invSboxRom_76;
      8'b01001101 : _zz_invSub_7 = invSboxRom_77;
      8'b01001110 : _zz_invSub_7 = invSboxRom_78;
      8'b01001111 : _zz_invSub_7 = invSboxRom_79;
      8'b01010000 : _zz_invSub_7 = invSboxRom_80;
      8'b01010001 : _zz_invSub_7 = invSboxRom_81;
      8'b01010010 : _zz_invSub_7 = invSboxRom_82;
      8'b01010011 : _zz_invSub_7 = invSboxRom_83;
      8'b01010100 : _zz_invSub_7 = invSboxRom_84;
      8'b01010101 : _zz_invSub_7 = invSboxRom_85;
      8'b01010110 : _zz_invSub_7 = invSboxRom_86;
      8'b01010111 : _zz_invSub_7 = invSboxRom_87;
      8'b01011000 : _zz_invSub_7 = invSboxRom_88;
      8'b01011001 : _zz_invSub_7 = invSboxRom_89;
      8'b01011010 : _zz_invSub_7 = invSboxRom_90;
      8'b01011011 : _zz_invSub_7 = invSboxRom_91;
      8'b01011100 : _zz_invSub_7 = invSboxRom_92;
      8'b01011101 : _zz_invSub_7 = invSboxRom_93;
      8'b01011110 : _zz_invSub_7 = invSboxRom_94;
      8'b01011111 : _zz_invSub_7 = invSboxRom_95;
      8'b01100000 : _zz_invSub_7 = invSboxRom_96;
      8'b01100001 : _zz_invSub_7 = invSboxRom_97;
      8'b01100010 : _zz_invSub_7 = invSboxRom_98;
      8'b01100011 : _zz_invSub_7 = invSboxRom_99;
      8'b01100100 : _zz_invSub_7 = invSboxRom_100;
      8'b01100101 : _zz_invSub_7 = invSboxRom_101;
      8'b01100110 : _zz_invSub_7 = invSboxRom_102;
      8'b01100111 : _zz_invSub_7 = invSboxRom_103;
      8'b01101000 : _zz_invSub_7 = invSboxRom_104;
      8'b01101001 : _zz_invSub_7 = invSboxRom_105;
      8'b01101010 : _zz_invSub_7 = invSboxRom_106;
      8'b01101011 : _zz_invSub_7 = invSboxRom_107;
      8'b01101100 : _zz_invSub_7 = invSboxRom_108;
      8'b01101101 : _zz_invSub_7 = invSboxRom_109;
      8'b01101110 : _zz_invSub_7 = invSboxRom_110;
      8'b01101111 : _zz_invSub_7 = invSboxRom_111;
      8'b01110000 : _zz_invSub_7 = invSboxRom_112;
      8'b01110001 : _zz_invSub_7 = invSboxRom_113;
      8'b01110010 : _zz_invSub_7 = invSboxRom_114;
      8'b01110011 : _zz_invSub_7 = invSboxRom_115;
      8'b01110100 : _zz_invSub_7 = invSboxRom_116;
      8'b01110101 : _zz_invSub_7 = invSboxRom_117;
      8'b01110110 : _zz_invSub_7 = invSboxRom_118;
      8'b01110111 : _zz_invSub_7 = invSboxRom_119;
      8'b01111000 : _zz_invSub_7 = invSboxRom_120;
      8'b01111001 : _zz_invSub_7 = invSboxRom_121;
      8'b01111010 : _zz_invSub_7 = invSboxRom_122;
      8'b01111011 : _zz_invSub_7 = invSboxRom_123;
      8'b01111100 : _zz_invSub_7 = invSboxRom_124;
      8'b01111101 : _zz_invSub_7 = invSboxRom_125;
      8'b01111110 : _zz_invSub_7 = invSboxRom_126;
      8'b01111111 : _zz_invSub_7 = invSboxRom_127;
      8'b10000000 : _zz_invSub_7 = invSboxRom_128;
      8'b10000001 : _zz_invSub_7 = invSboxRom_129;
      8'b10000010 : _zz_invSub_7 = invSboxRom_130;
      8'b10000011 : _zz_invSub_7 = invSboxRom_131;
      8'b10000100 : _zz_invSub_7 = invSboxRom_132;
      8'b10000101 : _zz_invSub_7 = invSboxRom_133;
      8'b10000110 : _zz_invSub_7 = invSboxRom_134;
      8'b10000111 : _zz_invSub_7 = invSboxRom_135;
      8'b10001000 : _zz_invSub_7 = invSboxRom_136;
      8'b10001001 : _zz_invSub_7 = invSboxRom_137;
      8'b10001010 : _zz_invSub_7 = invSboxRom_138;
      8'b10001011 : _zz_invSub_7 = invSboxRom_139;
      8'b10001100 : _zz_invSub_7 = invSboxRom_140;
      8'b10001101 : _zz_invSub_7 = invSboxRom_141;
      8'b10001110 : _zz_invSub_7 = invSboxRom_142;
      8'b10001111 : _zz_invSub_7 = invSboxRom_143;
      8'b10010000 : _zz_invSub_7 = invSboxRom_144;
      8'b10010001 : _zz_invSub_7 = invSboxRom_145;
      8'b10010010 : _zz_invSub_7 = invSboxRom_146;
      8'b10010011 : _zz_invSub_7 = invSboxRom_147;
      8'b10010100 : _zz_invSub_7 = invSboxRom_148;
      8'b10010101 : _zz_invSub_7 = invSboxRom_149;
      8'b10010110 : _zz_invSub_7 = invSboxRom_150;
      8'b10010111 : _zz_invSub_7 = invSboxRom_151;
      8'b10011000 : _zz_invSub_7 = invSboxRom_152;
      8'b10011001 : _zz_invSub_7 = invSboxRom_153;
      8'b10011010 : _zz_invSub_7 = invSboxRom_154;
      8'b10011011 : _zz_invSub_7 = invSboxRom_155;
      8'b10011100 : _zz_invSub_7 = invSboxRom_156;
      8'b10011101 : _zz_invSub_7 = invSboxRom_157;
      8'b10011110 : _zz_invSub_7 = invSboxRom_158;
      8'b10011111 : _zz_invSub_7 = invSboxRom_159;
      8'b10100000 : _zz_invSub_7 = invSboxRom_160;
      8'b10100001 : _zz_invSub_7 = invSboxRom_161;
      8'b10100010 : _zz_invSub_7 = invSboxRom_162;
      8'b10100011 : _zz_invSub_7 = invSboxRom_163;
      8'b10100100 : _zz_invSub_7 = invSboxRom_164;
      8'b10100101 : _zz_invSub_7 = invSboxRom_165;
      8'b10100110 : _zz_invSub_7 = invSboxRom_166;
      8'b10100111 : _zz_invSub_7 = invSboxRom_167;
      8'b10101000 : _zz_invSub_7 = invSboxRom_168;
      8'b10101001 : _zz_invSub_7 = invSboxRom_169;
      8'b10101010 : _zz_invSub_7 = invSboxRom_170;
      8'b10101011 : _zz_invSub_7 = invSboxRom_171;
      8'b10101100 : _zz_invSub_7 = invSboxRom_172;
      8'b10101101 : _zz_invSub_7 = invSboxRom_173;
      8'b10101110 : _zz_invSub_7 = invSboxRom_174;
      8'b10101111 : _zz_invSub_7 = invSboxRom_175;
      8'b10110000 : _zz_invSub_7 = invSboxRom_176;
      8'b10110001 : _zz_invSub_7 = invSboxRom_177;
      8'b10110010 : _zz_invSub_7 = invSboxRom_178;
      8'b10110011 : _zz_invSub_7 = invSboxRom_179;
      8'b10110100 : _zz_invSub_7 = invSboxRom_180;
      8'b10110101 : _zz_invSub_7 = invSboxRom_181;
      8'b10110110 : _zz_invSub_7 = invSboxRom_182;
      8'b10110111 : _zz_invSub_7 = invSboxRom_183;
      8'b10111000 : _zz_invSub_7 = invSboxRom_184;
      8'b10111001 : _zz_invSub_7 = invSboxRom_185;
      8'b10111010 : _zz_invSub_7 = invSboxRom_186;
      8'b10111011 : _zz_invSub_7 = invSboxRom_187;
      8'b10111100 : _zz_invSub_7 = invSboxRom_188;
      8'b10111101 : _zz_invSub_7 = invSboxRom_189;
      8'b10111110 : _zz_invSub_7 = invSboxRom_190;
      8'b10111111 : _zz_invSub_7 = invSboxRom_191;
      8'b11000000 : _zz_invSub_7 = invSboxRom_192;
      8'b11000001 : _zz_invSub_7 = invSboxRom_193;
      8'b11000010 : _zz_invSub_7 = invSboxRom_194;
      8'b11000011 : _zz_invSub_7 = invSboxRom_195;
      8'b11000100 : _zz_invSub_7 = invSboxRom_196;
      8'b11000101 : _zz_invSub_7 = invSboxRom_197;
      8'b11000110 : _zz_invSub_7 = invSboxRom_198;
      8'b11000111 : _zz_invSub_7 = invSboxRom_199;
      8'b11001000 : _zz_invSub_7 = invSboxRom_200;
      8'b11001001 : _zz_invSub_7 = invSboxRom_201;
      8'b11001010 : _zz_invSub_7 = invSboxRom_202;
      8'b11001011 : _zz_invSub_7 = invSboxRom_203;
      8'b11001100 : _zz_invSub_7 = invSboxRom_204;
      8'b11001101 : _zz_invSub_7 = invSboxRom_205;
      8'b11001110 : _zz_invSub_7 = invSboxRom_206;
      8'b11001111 : _zz_invSub_7 = invSboxRom_207;
      8'b11010000 : _zz_invSub_7 = invSboxRom_208;
      8'b11010001 : _zz_invSub_7 = invSboxRom_209;
      8'b11010010 : _zz_invSub_7 = invSboxRom_210;
      8'b11010011 : _zz_invSub_7 = invSboxRom_211;
      8'b11010100 : _zz_invSub_7 = invSboxRom_212;
      8'b11010101 : _zz_invSub_7 = invSboxRom_213;
      8'b11010110 : _zz_invSub_7 = invSboxRom_214;
      8'b11010111 : _zz_invSub_7 = invSboxRom_215;
      8'b11011000 : _zz_invSub_7 = invSboxRom_216;
      8'b11011001 : _zz_invSub_7 = invSboxRom_217;
      8'b11011010 : _zz_invSub_7 = invSboxRom_218;
      8'b11011011 : _zz_invSub_7 = invSboxRom_219;
      8'b11011100 : _zz_invSub_7 = invSboxRom_220;
      8'b11011101 : _zz_invSub_7 = invSboxRom_221;
      8'b11011110 : _zz_invSub_7 = invSboxRom_222;
      8'b11011111 : _zz_invSub_7 = invSboxRom_223;
      8'b11100000 : _zz_invSub_7 = invSboxRom_224;
      8'b11100001 : _zz_invSub_7 = invSboxRom_225;
      8'b11100010 : _zz_invSub_7 = invSboxRom_226;
      8'b11100011 : _zz_invSub_7 = invSboxRom_227;
      8'b11100100 : _zz_invSub_7 = invSboxRom_228;
      8'b11100101 : _zz_invSub_7 = invSboxRom_229;
      8'b11100110 : _zz_invSub_7 = invSboxRom_230;
      8'b11100111 : _zz_invSub_7 = invSboxRom_231;
      8'b11101000 : _zz_invSub_7 = invSboxRom_232;
      8'b11101001 : _zz_invSub_7 = invSboxRom_233;
      8'b11101010 : _zz_invSub_7 = invSboxRom_234;
      8'b11101011 : _zz_invSub_7 = invSboxRom_235;
      8'b11101100 : _zz_invSub_7 = invSboxRom_236;
      8'b11101101 : _zz_invSub_7 = invSboxRom_237;
      8'b11101110 : _zz_invSub_7 = invSboxRom_238;
      8'b11101111 : _zz_invSub_7 = invSboxRom_239;
      8'b11110000 : _zz_invSub_7 = invSboxRom_240;
      8'b11110001 : _zz_invSub_7 = invSboxRom_241;
      8'b11110010 : _zz_invSub_7 = invSboxRom_242;
      8'b11110011 : _zz_invSub_7 = invSboxRom_243;
      8'b11110100 : _zz_invSub_7 = invSboxRom_244;
      8'b11110101 : _zz_invSub_7 = invSboxRom_245;
      8'b11110110 : _zz_invSub_7 = invSboxRom_246;
      8'b11110111 : _zz_invSub_7 = invSboxRom_247;
      8'b11111000 : _zz_invSub_7 = invSboxRom_248;
      8'b11111001 : _zz_invSub_7 = invSboxRom_249;
      8'b11111010 : _zz_invSub_7 = invSboxRom_250;
      8'b11111011 : _zz_invSub_7 = invSboxRom_251;
      8'b11111100 : _zz_invSub_7 = invSboxRom_252;
      8'b11111101 : _zz_invSub_7 = invSboxRom_253;
      8'b11111110 : _zz_invSub_7 = invSboxRom_254;
      default : _zz_invSub_7 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_8)
      8'b00000000 : _zz_invSub_8 = invSboxRom_0;
      8'b00000001 : _zz_invSub_8 = invSboxRom_1;
      8'b00000010 : _zz_invSub_8 = invSboxRom_2;
      8'b00000011 : _zz_invSub_8 = invSboxRom_3;
      8'b00000100 : _zz_invSub_8 = invSboxRom_4;
      8'b00000101 : _zz_invSub_8 = invSboxRom_5;
      8'b00000110 : _zz_invSub_8 = invSboxRom_6;
      8'b00000111 : _zz_invSub_8 = invSboxRom_7;
      8'b00001000 : _zz_invSub_8 = invSboxRom_8;
      8'b00001001 : _zz_invSub_8 = invSboxRom_9;
      8'b00001010 : _zz_invSub_8 = invSboxRom_10;
      8'b00001011 : _zz_invSub_8 = invSboxRom_11;
      8'b00001100 : _zz_invSub_8 = invSboxRom_12;
      8'b00001101 : _zz_invSub_8 = invSboxRom_13;
      8'b00001110 : _zz_invSub_8 = invSboxRom_14;
      8'b00001111 : _zz_invSub_8 = invSboxRom_15;
      8'b00010000 : _zz_invSub_8 = invSboxRom_16;
      8'b00010001 : _zz_invSub_8 = invSboxRom_17;
      8'b00010010 : _zz_invSub_8 = invSboxRom_18;
      8'b00010011 : _zz_invSub_8 = invSboxRom_19;
      8'b00010100 : _zz_invSub_8 = invSboxRom_20;
      8'b00010101 : _zz_invSub_8 = invSboxRom_21;
      8'b00010110 : _zz_invSub_8 = invSboxRom_22;
      8'b00010111 : _zz_invSub_8 = invSboxRom_23;
      8'b00011000 : _zz_invSub_8 = invSboxRom_24;
      8'b00011001 : _zz_invSub_8 = invSboxRom_25;
      8'b00011010 : _zz_invSub_8 = invSboxRom_26;
      8'b00011011 : _zz_invSub_8 = invSboxRom_27;
      8'b00011100 : _zz_invSub_8 = invSboxRom_28;
      8'b00011101 : _zz_invSub_8 = invSboxRom_29;
      8'b00011110 : _zz_invSub_8 = invSboxRom_30;
      8'b00011111 : _zz_invSub_8 = invSboxRom_31;
      8'b00100000 : _zz_invSub_8 = invSboxRom_32;
      8'b00100001 : _zz_invSub_8 = invSboxRom_33;
      8'b00100010 : _zz_invSub_8 = invSboxRom_34;
      8'b00100011 : _zz_invSub_8 = invSboxRom_35;
      8'b00100100 : _zz_invSub_8 = invSboxRom_36;
      8'b00100101 : _zz_invSub_8 = invSboxRom_37;
      8'b00100110 : _zz_invSub_8 = invSboxRom_38;
      8'b00100111 : _zz_invSub_8 = invSboxRom_39;
      8'b00101000 : _zz_invSub_8 = invSboxRom_40;
      8'b00101001 : _zz_invSub_8 = invSboxRom_41;
      8'b00101010 : _zz_invSub_8 = invSboxRom_42;
      8'b00101011 : _zz_invSub_8 = invSboxRom_43;
      8'b00101100 : _zz_invSub_8 = invSboxRom_44;
      8'b00101101 : _zz_invSub_8 = invSboxRom_45;
      8'b00101110 : _zz_invSub_8 = invSboxRom_46;
      8'b00101111 : _zz_invSub_8 = invSboxRom_47;
      8'b00110000 : _zz_invSub_8 = invSboxRom_48;
      8'b00110001 : _zz_invSub_8 = invSboxRom_49;
      8'b00110010 : _zz_invSub_8 = invSboxRom_50;
      8'b00110011 : _zz_invSub_8 = invSboxRom_51;
      8'b00110100 : _zz_invSub_8 = invSboxRom_52;
      8'b00110101 : _zz_invSub_8 = invSboxRom_53;
      8'b00110110 : _zz_invSub_8 = invSboxRom_54;
      8'b00110111 : _zz_invSub_8 = invSboxRom_55;
      8'b00111000 : _zz_invSub_8 = invSboxRom_56;
      8'b00111001 : _zz_invSub_8 = invSboxRom_57;
      8'b00111010 : _zz_invSub_8 = invSboxRom_58;
      8'b00111011 : _zz_invSub_8 = invSboxRom_59;
      8'b00111100 : _zz_invSub_8 = invSboxRom_60;
      8'b00111101 : _zz_invSub_8 = invSboxRom_61;
      8'b00111110 : _zz_invSub_8 = invSboxRom_62;
      8'b00111111 : _zz_invSub_8 = invSboxRom_63;
      8'b01000000 : _zz_invSub_8 = invSboxRom_64;
      8'b01000001 : _zz_invSub_8 = invSboxRom_65;
      8'b01000010 : _zz_invSub_8 = invSboxRom_66;
      8'b01000011 : _zz_invSub_8 = invSboxRom_67;
      8'b01000100 : _zz_invSub_8 = invSboxRom_68;
      8'b01000101 : _zz_invSub_8 = invSboxRom_69;
      8'b01000110 : _zz_invSub_8 = invSboxRom_70;
      8'b01000111 : _zz_invSub_8 = invSboxRom_71;
      8'b01001000 : _zz_invSub_8 = invSboxRom_72;
      8'b01001001 : _zz_invSub_8 = invSboxRom_73;
      8'b01001010 : _zz_invSub_8 = invSboxRom_74;
      8'b01001011 : _zz_invSub_8 = invSboxRom_75;
      8'b01001100 : _zz_invSub_8 = invSboxRom_76;
      8'b01001101 : _zz_invSub_8 = invSboxRom_77;
      8'b01001110 : _zz_invSub_8 = invSboxRom_78;
      8'b01001111 : _zz_invSub_8 = invSboxRom_79;
      8'b01010000 : _zz_invSub_8 = invSboxRom_80;
      8'b01010001 : _zz_invSub_8 = invSboxRom_81;
      8'b01010010 : _zz_invSub_8 = invSboxRom_82;
      8'b01010011 : _zz_invSub_8 = invSboxRom_83;
      8'b01010100 : _zz_invSub_8 = invSboxRom_84;
      8'b01010101 : _zz_invSub_8 = invSboxRom_85;
      8'b01010110 : _zz_invSub_8 = invSboxRom_86;
      8'b01010111 : _zz_invSub_8 = invSboxRom_87;
      8'b01011000 : _zz_invSub_8 = invSboxRom_88;
      8'b01011001 : _zz_invSub_8 = invSboxRom_89;
      8'b01011010 : _zz_invSub_8 = invSboxRom_90;
      8'b01011011 : _zz_invSub_8 = invSboxRom_91;
      8'b01011100 : _zz_invSub_8 = invSboxRom_92;
      8'b01011101 : _zz_invSub_8 = invSboxRom_93;
      8'b01011110 : _zz_invSub_8 = invSboxRom_94;
      8'b01011111 : _zz_invSub_8 = invSboxRom_95;
      8'b01100000 : _zz_invSub_8 = invSboxRom_96;
      8'b01100001 : _zz_invSub_8 = invSboxRom_97;
      8'b01100010 : _zz_invSub_8 = invSboxRom_98;
      8'b01100011 : _zz_invSub_8 = invSboxRom_99;
      8'b01100100 : _zz_invSub_8 = invSboxRom_100;
      8'b01100101 : _zz_invSub_8 = invSboxRom_101;
      8'b01100110 : _zz_invSub_8 = invSboxRom_102;
      8'b01100111 : _zz_invSub_8 = invSboxRom_103;
      8'b01101000 : _zz_invSub_8 = invSboxRom_104;
      8'b01101001 : _zz_invSub_8 = invSboxRom_105;
      8'b01101010 : _zz_invSub_8 = invSboxRom_106;
      8'b01101011 : _zz_invSub_8 = invSboxRom_107;
      8'b01101100 : _zz_invSub_8 = invSboxRom_108;
      8'b01101101 : _zz_invSub_8 = invSboxRom_109;
      8'b01101110 : _zz_invSub_8 = invSboxRom_110;
      8'b01101111 : _zz_invSub_8 = invSboxRom_111;
      8'b01110000 : _zz_invSub_8 = invSboxRom_112;
      8'b01110001 : _zz_invSub_8 = invSboxRom_113;
      8'b01110010 : _zz_invSub_8 = invSboxRom_114;
      8'b01110011 : _zz_invSub_8 = invSboxRom_115;
      8'b01110100 : _zz_invSub_8 = invSboxRom_116;
      8'b01110101 : _zz_invSub_8 = invSboxRom_117;
      8'b01110110 : _zz_invSub_8 = invSboxRom_118;
      8'b01110111 : _zz_invSub_8 = invSboxRom_119;
      8'b01111000 : _zz_invSub_8 = invSboxRom_120;
      8'b01111001 : _zz_invSub_8 = invSboxRom_121;
      8'b01111010 : _zz_invSub_8 = invSboxRom_122;
      8'b01111011 : _zz_invSub_8 = invSboxRom_123;
      8'b01111100 : _zz_invSub_8 = invSboxRom_124;
      8'b01111101 : _zz_invSub_8 = invSboxRom_125;
      8'b01111110 : _zz_invSub_8 = invSboxRom_126;
      8'b01111111 : _zz_invSub_8 = invSboxRom_127;
      8'b10000000 : _zz_invSub_8 = invSboxRom_128;
      8'b10000001 : _zz_invSub_8 = invSboxRom_129;
      8'b10000010 : _zz_invSub_8 = invSboxRom_130;
      8'b10000011 : _zz_invSub_8 = invSboxRom_131;
      8'b10000100 : _zz_invSub_8 = invSboxRom_132;
      8'b10000101 : _zz_invSub_8 = invSboxRom_133;
      8'b10000110 : _zz_invSub_8 = invSboxRom_134;
      8'b10000111 : _zz_invSub_8 = invSboxRom_135;
      8'b10001000 : _zz_invSub_8 = invSboxRom_136;
      8'b10001001 : _zz_invSub_8 = invSboxRom_137;
      8'b10001010 : _zz_invSub_8 = invSboxRom_138;
      8'b10001011 : _zz_invSub_8 = invSboxRom_139;
      8'b10001100 : _zz_invSub_8 = invSboxRom_140;
      8'b10001101 : _zz_invSub_8 = invSboxRom_141;
      8'b10001110 : _zz_invSub_8 = invSboxRom_142;
      8'b10001111 : _zz_invSub_8 = invSboxRom_143;
      8'b10010000 : _zz_invSub_8 = invSboxRom_144;
      8'b10010001 : _zz_invSub_8 = invSboxRom_145;
      8'b10010010 : _zz_invSub_8 = invSboxRom_146;
      8'b10010011 : _zz_invSub_8 = invSboxRom_147;
      8'b10010100 : _zz_invSub_8 = invSboxRom_148;
      8'b10010101 : _zz_invSub_8 = invSboxRom_149;
      8'b10010110 : _zz_invSub_8 = invSboxRom_150;
      8'b10010111 : _zz_invSub_8 = invSboxRom_151;
      8'b10011000 : _zz_invSub_8 = invSboxRom_152;
      8'b10011001 : _zz_invSub_8 = invSboxRom_153;
      8'b10011010 : _zz_invSub_8 = invSboxRom_154;
      8'b10011011 : _zz_invSub_8 = invSboxRom_155;
      8'b10011100 : _zz_invSub_8 = invSboxRom_156;
      8'b10011101 : _zz_invSub_8 = invSboxRom_157;
      8'b10011110 : _zz_invSub_8 = invSboxRom_158;
      8'b10011111 : _zz_invSub_8 = invSboxRom_159;
      8'b10100000 : _zz_invSub_8 = invSboxRom_160;
      8'b10100001 : _zz_invSub_8 = invSboxRom_161;
      8'b10100010 : _zz_invSub_8 = invSboxRom_162;
      8'b10100011 : _zz_invSub_8 = invSboxRom_163;
      8'b10100100 : _zz_invSub_8 = invSboxRom_164;
      8'b10100101 : _zz_invSub_8 = invSboxRom_165;
      8'b10100110 : _zz_invSub_8 = invSboxRom_166;
      8'b10100111 : _zz_invSub_8 = invSboxRom_167;
      8'b10101000 : _zz_invSub_8 = invSboxRom_168;
      8'b10101001 : _zz_invSub_8 = invSboxRom_169;
      8'b10101010 : _zz_invSub_8 = invSboxRom_170;
      8'b10101011 : _zz_invSub_8 = invSboxRom_171;
      8'b10101100 : _zz_invSub_8 = invSboxRom_172;
      8'b10101101 : _zz_invSub_8 = invSboxRom_173;
      8'b10101110 : _zz_invSub_8 = invSboxRom_174;
      8'b10101111 : _zz_invSub_8 = invSboxRom_175;
      8'b10110000 : _zz_invSub_8 = invSboxRom_176;
      8'b10110001 : _zz_invSub_8 = invSboxRom_177;
      8'b10110010 : _zz_invSub_8 = invSboxRom_178;
      8'b10110011 : _zz_invSub_8 = invSboxRom_179;
      8'b10110100 : _zz_invSub_8 = invSboxRom_180;
      8'b10110101 : _zz_invSub_8 = invSboxRom_181;
      8'b10110110 : _zz_invSub_8 = invSboxRom_182;
      8'b10110111 : _zz_invSub_8 = invSboxRom_183;
      8'b10111000 : _zz_invSub_8 = invSboxRom_184;
      8'b10111001 : _zz_invSub_8 = invSboxRom_185;
      8'b10111010 : _zz_invSub_8 = invSboxRom_186;
      8'b10111011 : _zz_invSub_8 = invSboxRom_187;
      8'b10111100 : _zz_invSub_8 = invSboxRom_188;
      8'b10111101 : _zz_invSub_8 = invSboxRom_189;
      8'b10111110 : _zz_invSub_8 = invSboxRom_190;
      8'b10111111 : _zz_invSub_8 = invSboxRom_191;
      8'b11000000 : _zz_invSub_8 = invSboxRom_192;
      8'b11000001 : _zz_invSub_8 = invSboxRom_193;
      8'b11000010 : _zz_invSub_8 = invSboxRom_194;
      8'b11000011 : _zz_invSub_8 = invSboxRom_195;
      8'b11000100 : _zz_invSub_8 = invSboxRom_196;
      8'b11000101 : _zz_invSub_8 = invSboxRom_197;
      8'b11000110 : _zz_invSub_8 = invSboxRom_198;
      8'b11000111 : _zz_invSub_8 = invSboxRom_199;
      8'b11001000 : _zz_invSub_8 = invSboxRom_200;
      8'b11001001 : _zz_invSub_8 = invSboxRom_201;
      8'b11001010 : _zz_invSub_8 = invSboxRom_202;
      8'b11001011 : _zz_invSub_8 = invSboxRom_203;
      8'b11001100 : _zz_invSub_8 = invSboxRom_204;
      8'b11001101 : _zz_invSub_8 = invSboxRom_205;
      8'b11001110 : _zz_invSub_8 = invSboxRom_206;
      8'b11001111 : _zz_invSub_8 = invSboxRom_207;
      8'b11010000 : _zz_invSub_8 = invSboxRom_208;
      8'b11010001 : _zz_invSub_8 = invSboxRom_209;
      8'b11010010 : _zz_invSub_8 = invSboxRom_210;
      8'b11010011 : _zz_invSub_8 = invSboxRom_211;
      8'b11010100 : _zz_invSub_8 = invSboxRom_212;
      8'b11010101 : _zz_invSub_8 = invSboxRom_213;
      8'b11010110 : _zz_invSub_8 = invSboxRom_214;
      8'b11010111 : _zz_invSub_8 = invSboxRom_215;
      8'b11011000 : _zz_invSub_8 = invSboxRom_216;
      8'b11011001 : _zz_invSub_8 = invSboxRom_217;
      8'b11011010 : _zz_invSub_8 = invSboxRom_218;
      8'b11011011 : _zz_invSub_8 = invSboxRom_219;
      8'b11011100 : _zz_invSub_8 = invSboxRom_220;
      8'b11011101 : _zz_invSub_8 = invSboxRom_221;
      8'b11011110 : _zz_invSub_8 = invSboxRom_222;
      8'b11011111 : _zz_invSub_8 = invSboxRom_223;
      8'b11100000 : _zz_invSub_8 = invSboxRom_224;
      8'b11100001 : _zz_invSub_8 = invSboxRom_225;
      8'b11100010 : _zz_invSub_8 = invSboxRom_226;
      8'b11100011 : _zz_invSub_8 = invSboxRom_227;
      8'b11100100 : _zz_invSub_8 = invSboxRom_228;
      8'b11100101 : _zz_invSub_8 = invSboxRom_229;
      8'b11100110 : _zz_invSub_8 = invSboxRom_230;
      8'b11100111 : _zz_invSub_8 = invSboxRom_231;
      8'b11101000 : _zz_invSub_8 = invSboxRom_232;
      8'b11101001 : _zz_invSub_8 = invSboxRom_233;
      8'b11101010 : _zz_invSub_8 = invSboxRom_234;
      8'b11101011 : _zz_invSub_8 = invSboxRom_235;
      8'b11101100 : _zz_invSub_8 = invSboxRom_236;
      8'b11101101 : _zz_invSub_8 = invSboxRom_237;
      8'b11101110 : _zz_invSub_8 = invSboxRom_238;
      8'b11101111 : _zz_invSub_8 = invSboxRom_239;
      8'b11110000 : _zz_invSub_8 = invSboxRom_240;
      8'b11110001 : _zz_invSub_8 = invSboxRom_241;
      8'b11110010 : _zz_invSub_8 = invSboxRom_242;
      8'b11110011 : _zz_invSub_8 = invSboxRom_243;
      8'b11110100 : _zz_invSub_8 = invSboxRom_244;
      8'b11110101 : _zz_invSub_8 = invSboxRom_245;
      8'b11110110 : _zz_invSub_8 = invSboxRom_246;
      8'b11110111 : _zz_invSub_8 = invSboxRom_247;
      8'b11111000 : _zz_invSub_8 = invSboxRom_248;
      8'b11111001 : _zz_invSub_8 = invSboxRom_249;
      8'b11111010 : _zz_invSub_8 = invSboxRom_250;
      8'b11111011 : _zz_invSub_8 = invSboxRom_251;
      8'b11111100 : _zz_invSub_8 = invSboxRom_252;
      8'b11111101 : _zz_invSub_8 = invSboxRom_253;
      8'b11111110 : _zz_invSub_8 = invSboxRom_254;
      default : _zz_invSub_8 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_9)
      8'b00000000 : _zz_invSub_9 = invSboxRom_0;
      8'b00000001 : _zz_invSub_9 = invSboxRom_1;
      8'b00000010 : _zz_invSub_9 = invSboxRom_2;
      8'b00000011 : _zz_invSub_9 = invSboxRom_3;
      8'b00000100 : _zz_invSub_9 = invSboxRom_4;
      8'b00000101 : _zz_invSub_9 = invSboxRom_5;
      8'b00000110 : _zz_invSub_9 = invSboxRom_6;
      8'b00000111 : _zz_invSub_9 = invSboxRom_7;
      8'b00001000 : _zz_invSub_9 = invSboxRom_8;
      8'b00001001 : _zz_invSub_9 = invSboxRom_9;
      8'b00001010 : _zz_invSub_9 = invSboxRom_10;
      8'b00001011 : _zz_invSub_9 = invSboxRom_11;
      8'b00001100 : _zz_invSub_9 = invSboxRom_12;
      8'b00001101 : _zz_invSub_9 = invSboxRom_13;
      8'b00001110 : _zz_invSub_9 = invSboxRom_14;
      8'b00001111 : _zz_invSub_9 = invSboxRom_15;
      8'b00010000 : _zz_invSub_9 = invSboxRom_16;
      8'b00010001 : _zz_invSub_9 = invSboxRom_17;
      8'b00010010 : _zz_invSub_9 = invSboxRom_18;
      8'b00010011 : _zz_invSub_9 = invSboxRom_19;
      8'b00010100 : _zz_invSub_9 = invSboxRom_20;
      8'b00010101 : _zz_invSub_9 = invSboxRom_21;
      8'b00010110 : _zz_invSub_9 = invSboxRom_22;
      8'b00010111 : _zz_invSub_9 = invSboxRom_23;
      8'b00011000 : _zz_invSub_9 = invSboxRom_24;
      8'b00011001 : _zz_invSub_9 = invSboxRom_25;
      8'b00011010 : _zz_invSub_9 = invSboxRom_26;
      8'b00011011 : _zz_invSub_9 = invSboxRom_27;
      8'b00011100 : _zz_invSub_9 = invSboxRom_28;
      8'b00011101 : _zz_invSub_9 = invSboxRom_29;
      8'b00011110 : _zz_invSub_9 = invSboxRom_30;
      8'b00011111 : _zz_invSub_9 = invSboxRom_31;
      8'b00100000 : _zz_invSub_9 = invSboxRom_32;
      8'b00100001 : _zz_invSub_9 = invSboxRom_33;
      8'b00100010 : _zz_invSub_9 = invSboxRom_34;
      8'b00100011 : _zz_invSub_9 = invSboxRom_35;
      8'b00100100 : _zz_invSub_9 = invSboxRom_36;
      8'b00100101 : _zz_invSub_9 = invSboxRom_37;
      8'b00100110 : _zz_invSub_9 = invSboxRom_38;
      8'b00100111 : _zz_invSub_9 = invSboxRom_39;
      8'b00101000 : _zz_invSub_9 = invSboxRom_40;
      8'b00101001 : _zz_invSub_9 = invSboxRom_41;
      8'b00101010 : _zz_invSub_9 = invSboxRom_42;
      8'b00101011 : _zz_invSub_9 = invSboxRom_43;
      8'b00101100 : _zz_invSub_9 = invSboxRom_44;
      8'b00101101 : _zz_invSub_9 = invSboxRom_45;
      8'b00101110 : _zz_invSub_9 = invSboxRom_46;
      8'b00101111 : _zz_invSub_9 = invSboxRom_47;
      8'b00110000 : _zz_invSub_9 = invSboxRom_48;
      8'b00110001 : _zz_invSub_9 = invSboxRom_49;
      8'b00110010 : _zz_invSub_9 = invSboxRom_50;
      8'b00110011 : _zz_invSub_9 = invSboxRom_51;
      8'b00110100 : _zz_invSub_9 = invSboxRom_52;
      8'b00110101 : _zz_invSub_9 = invSboxRom_53;
      8'b00110110 : _zz_invSub_9 = invSboxRom_54;
      8'b00110111 : _zz_invSub_9 = invSboxRom_55;
      8'b00111000 : _zz_invSub_9 = invSboxRom_56;
      8'b00111001 : _zz_invSub_9 = invSboxRom_57;
      8'b00111010 : _zz_invSub_9 = invSboxRom_58;
      8'b00111011 : _zz_invSub_9 = invSboxRom_59;
      8'b00111100 : _zz_invSub_9 = invSboxRom_60;
      8'b00111101 : _zz_invSub_9 = invSboxRom_61;
      8'b00111110 : _zz_invSub_9 = invSboxRom_62;
      8'b00111111 : _zz_invSub_9 = invSboxRom_63;
      8'b01000000 : _zz_invSub_9 = invSboxRom_64;
      8'b01000001 : _zz_invSub_9 = invSboxRom_65;
      8'b01000010 : _zz_invSub_9 = invSboxRom_66;
      8'b01000011 : _zz_invSub_9 = invSboxRom_67;
      8'b01000100 : _zz_invSub_9 = invSboxRom_68;
      8'b01000101 : _zz_invSub_9 = invSboxRom_69;
      8'b01000110 : _zz_invSub_9 = invSboxRom_70;
      8'b01000111 : _zz_invSub_9 = invSboxRom_71;
      8'b01001000 : _zz_invSub_9 = invSboxRom_72;
      8'b01001001 : _zz_invSub_9 = invSboxRom_73;
      8'b01001010 : _zz_invSub_9 = invSboxRom_74;
      8'b01001011 : _zz_invSub_9 = invSboxRom_75;
      8'b01001100 : _zz_invSub_9 = invSboxRom_76;
      8'b01001101 : _zz_invSub_9 = invSboxRom_77;
      8'b01001110 : _zz_invSub_9 = invSboxRom_78;
      8'b01001111 : _zz_invSub_9 = invSboxRom_79;
      8'b01010000 : _zz_invSub_9 = invSboxRom_80;
      8'b01010001 : _zz_invSub_9 = invSboxRom_81;
      8'b01010010 : _zz_invSub_9 = invSboxRom_82;
      8'b01010011 : _zz_invSub_9 = invSboxRom_83;
      8'b01010100 : _zz_invSub_9 = invSboxRom_84;
      8'b01010101 : _zz_invSub_9 = invSboxRom_85;
      8'b01010110 : _zz_invSub_9 = invSboxRom_86;
      8'b01010111 : _zz_invSub_9 = invSboxRom_87;
      8'b01011000 : _zz_invSub_9 = invSboxRom_88;
      8'b01011001 : _zz_invSub_9 = invSboxRom_89;
      8'b01011010 : _zz_invSub_9 = invSboxRom_90;
      8'b01011011 : _zz_invSub_9 = invSboxRom_91;
      8'b01011100 : _zz_invSub_9 = invSboxRom_92;
      8'b01011101 : _zz_invSub_9 = invSboxRom_93;
      8'b01011110 : _zz_invSub_9 = invSboxRom_94;
      8'b01011111 : _zz_invSub_9 = invSboxRom_95;
      8'b01100000 : _zz_invSub_9 = invSboxRom_96;
      8'b01100001 : _zz_invSub_9 = invSboxRom_97;
      8'b01100010 : _zz_invSub_9 = invSboxRom_98;
      8'b01100011 : _zz_invSub_9 = invSboxRom_99;
      8'b01100100 : _zz_invSub_9 = invSboxRom_100;
      8'b01100101 : _zz_invSub_9 = invSboxRom_101;
      8'b01100110 : _zz_invSub_9 = invSboxRom_102;
      8'b01100111 : _zz_invSub_9 = invSboxRom_103;
      8'b01101000 : _zz_invSub_9 = invSboxRom_104;
      8'b01101001 : _zz_invSub_9 = invSboxRom_105;
      8'b01101010 : _zz_invSub_9 = invSboxRom_106;
      8'b01101011 : _zz_invSub_9 = invSboxRom_107;
      8'b01101100 : _zz_invSub_9 = invSboxRom_108;
      8'b01101101 : _zz_invSub_9 = invSboxRom_109;
      8'b01101110 : _zz_invSub_9 = invSboxRom_110;
      8'b01101111 : _zz_invSub_9 = invSboxRom_111;
      8'b01110000 : _zz_invSub_9 = invSboxRom_112;
      8'b01110001 : _zz_invSub_9 = invSboxRom_113;
      8'b01110010 : _zz_invSub_9 = invSboxRom_114;
      8'b01110011 : _zz_invSub_9 = invSboxRom_115;
      8'b01110100 : _zz_invSub_9 = invSboxRom_116;
      8'b01110101 : _zz_invSub_9 = invSboxRom_117;
      8'b01110110 : _zz_invSub_9 = invSboxRom_118;
      8'b01110111 : _zz_invSub_9 = invSboxRom_119;
      8'b01111000 : _zz_invSub_9 = invSboxRom_120;
      8'b01111001 : _zz_invSub_9 = invSboxRom_121;
      8'b01111010 : _zz_invSub_9 = invSboxRom_122;
      8'b01111011 : _zz_invSub_9 = invSboxRom_123;
      8'b01111100 : _zz_invSub_9 = invSboxRom_124;
      8'b01111101 : _zz_invSub_9 = invSboxRom_125;
      8'b01111110 : _zz_invSub_9 = invSboxRom_126;
      8'b01111111 : _zz_invSub_9 = invSboxRom_127;
      8'b10000000 : _zz_invSub_9 = invSboxRom_128;
      8'b10000001 : _zz_invSub_9 = invSboxRom_129;
      8'b10000010 : _zz_invSub_9 = invSboxRom_130;
      8'b10000011 : _zz_invSub_9 = invSboxRom_131;
      8'b10000100 : _zz_invSub_9 = invSboxRom_132;
      8'b10000101 : _zz_invSub_9 = invSboxRom_133;
      8'b10000110 : _zz_invSub_9 = invSboxRom_134;
      8'b10000111 : _zz_invSub_9 = invSboxRom_135;
      8'b10001000 : _zz_invSub_9 = invSboxRom_136;
      8'b10001001 : _zz_invSub_9 = invSboxRom_137;
      8'b10001010 : _zz_invSub_9 = invSboxRom_138;
      8'b10001011 : _zz_invSub_9 = invSboxRom_139;
      8'b10001100 : _zz_invSub_9 = invSboxRom_140;
      8'b10001101 : _zz_invSub_9 = invSboxRom_141;
      8'b10001110 : _zz_invSub_9 = invSboxRom_142;
      8'b10001111 : _zz_invSub_9 = invSboxRom_143;
      8'b10010000 : _zz_invSub_9 = invSboxRom_144;
      8'b10010001 : _zz_invSub_9 = invSboxRom_145;
      8'b10010010 : _zz_invSub_9 = invSboxRom_146;
      8'b10010011 : _zz_invSub_9 = invSboxRom_147;
      8'b10010100 : _zz_invSub_9 = invSboxRom_148;
      8'b10010101 : _zz_invSub_9 = invSboxRom_149;
      8'b10010110 : _zz_invSub_9 = invSboxRom_150;
      8'b10010111 : _zz_invSub_9 = invSboxRom_151;
      8'b10011000 : _zz_invSub_9 = invSboxRom_152;
      8'b10011001 : _zz_invSub_9 = invSboxRom_153;
      8'b10011010 : _zz_invSub_9 = invSboxRom_154;
      8'b10011011 : _zz_invSub_9 = invSboxRom_155;
      8'b10011100 : _zz_invSub_9 = invSboxRom_156;
      8'b10011101 : _zz_invSub_9 = invSboxRom_157;
      8'b10011110 : _zz_invSub_9 = invSboxRom_158;
      8'b10011111 : _zz_invSub_9 = invSboxRom_159;
      8'b10100000 : _zz_invSub_9 = invSboxRom_160;
      8'b10100001 : _zz_invSub_9 = invSboxRom_161;
      8'b10100010 : _zz_invSub_9 = invSboxRom_162;
      8'b10100011 : _zz_invSub_9 = invSboxRom_163;
      8'b10100100 : _zz_invSub_9 = invSboxRom_164;
      8'b10100101 : _zz_invSub_9 = invSboxRom_165;
      8'b10100110 : _zz_invSub_9 = invSboxRom_166;
      8'b10100111 : _zz_invSub_9 = invSboxRom_167;
      8'b10101000 : _zz_invSub_9 = invSboxRom_168;
      8'b10101001 : _zz_invSub_9 = invSboxRom_169;
      8'b10101010 : _zz_invSub_9 = invSboxRom_170;
      8'b10101011 : _zz_invSub_9 = invSboxRom_171;
      8'b10101100 : _zz_invSub_9 = invSboxRom_172;
      8'b10101101 : _zz_invSub_9 = invSboxRom_173;
      8'b10101110 : _zz_invSub_9 = invSboxRom_174;
      8'b10101111 : _zz_invSub_9 = invSboxRom_175;
      8'b10110000 : _zz_invSub_9 = invSboxRom_176;
      8'b10110001 : _zz_invSub_9 = invSboxRom_177;
      8'b10110010 : _zz_invSub_9 = invSboxRom_178;
      8'b10110011 : _zz_invSub_9 = invSboxRom_179;
      8'b10110100 : _zz_invSub_9 = invSboxRom_180;
      8'b10110101 : _zz_invSub_9 = invSboxRom_181;
      8'b10110110 : _zz_invSub_9 = invSboxRom_182;
      8'b10110111 : _zz_invSub_9 = invSboxRom_183;
      8'b10111000 : _zz_invSub_9 = invSboxRom_184;
      8'b10111001 : _zz_invSub_9 = invSboxRom_185;
      8'b10111010 : _zz_invSub_9 = invSboxRom_186;
      8'b10111011 : _zz_invSub_9 = invSboxRom_187;
      8'b10111100 : _zz_invSub_9 = invSboxRom_188;
      8'b10111101 : _zz_invSub_9 = invSboxRom_189;
      8'b10111110 : _zz_invSub_9 = invSboxRom_190;
      8'b10111111 : _zz_invSub_9 = invSboxRom_191;
      8'b11000000 : _zz_invSub_9 = invSboxRom_192;
      8'b11000001 : _zz_invSub_9 = invSboxRom_193;
      8'b11000010 : _zz_invSub_9 = invSboxRom_194;
      8'b11000011 : _zz_invSub_9 = invSboxRom_195;
      8'b11000100 : _zz_invSub_9 = invSboxRom_196;
      8'b11000101 : _zz_invSub_9 = invSboxRom_197;
      8'b11000110 : _zz_invSub_9 = invSboxRom_198;
      8'b11000111 : _zz_invSub_9 = invSboxRom_199;
      8'b11001000 : _zz_invSub_9 = invSboxRom_200;
      8'b11001001 : _zz_invSub_9 = invSboxRom_201;
      8'b11001010 : _zz_invSub_9 = invSboxRom_202;
      8'b11001011 : _zz_invSub_9 = invSboxRom_203;
      8'b11001100 : _zz_invSub_9 = invSboxRom_204;
      8'b11001101 : _zz_invSub_9 = invSboxRom_205;
      8'b11001110 : _zz_invSub_9 = invSboxRom_206;
      8'b11001111 : _zz_invSub_9 = invSboxRom_207;
      8'b11010000 : _zz_invSub_9 = invSboxRom_208;
      8'b11010001 : _zz_invSub_9 = invSboxRom_209;
      8'b11010010 : _zz_invSub_9 = invSboxRom_210;
      8'b11010011 : _zz_invSub_9 = invSboxRom_211;
      8'b11010100 : _zz_invSub_9 = invSboxRom_212;
      8'b11010101 : _zz_invSub_9 = invSboxRom_213;
      8'b11010110 : _zz_invSub_9 = invSboxRom_214;
      8'b11010111 : _zz_invSub_9 = invSboxRom_215;
      8'b11011000 : _zz_invSub_9 = invSboxRom_216;
      8'b11011001 : _zz_invSub_9 = invSboxRom_217;
      8'b11011010 : _zz_invSub_9 = invSboxRom_218;
      8'b11011011 : _zz_invSub_9 = invSboxRom_219;
      8'b11011100 : _zz_invSub_9 = invSboxRom_220;
      8'b11011101 : _zz_invSub_9 = invSboxRom_221;
      8'b11011110 : _zz_invSub_9 = invSboxRom_222;
      8'b11011111 : _zz_invSub_9 = invSboxRom_223;
      8'b11100000 : _zz_invSub_9 = invSboxRom_224;
      8'b11100001 : _zz_invSub_9 = invSboxRom_225;
      8'b11100010 : _zz_invSub_9 = invSboxRom_226;
      8'b11100011 : _zz_invSub_9 = invSboxRom_227;
      8'b11100100 : _zz_invSub_9 = invSboxRom_228;
      8'b11100101 : _zz_invSub_9 = invSboxRom_229;
      8'b11100110 : _zz_invSub_9 = invSboxRom_230;
      8'b11100111 : _zz_invSub_9 = invSboxRom_231;
      8'b11101000 : _zz_invSub_9 = invSboxRom_232;
      8'b11101001 : _zz_invSub_9 = invSboxRom_233;
      8'b11101010 : _zz_invSub_9 = invSboxRom_234;
      8'b11101011 : _zz_invSub_9 = invSboxRom_235;
      8'b11101100 : _zz_invSub_9 = invSboxRom_236;
      8'b11101101 : _zz_invSub_9 = invSboxRom_237;
      8'b11101110 : _zz_invSub_9 = invSboxRom_238;
      8'b11101111 : _zz_invSub_9 = invSboxRom_239;
      8'b11110000 : _zz_invSub_9 = invSboxRom_240;
      8'b11110001 : _zz_invSub_9 = invSboxRom_241;
      8'b11110010 : _zz_invSub_9 = invSboxRom_242;
      8'b11110011 : _zz_invSub_9 = invSboxRom_243;
      8'b11110100 : _zz_invSub_9 = invSboxRom_244;
      8'b11110101 : _zz_invSub_9 = invSboxRom_245;
      8'b11110110 : _zz_invSub_9 = invSboxRom_246;
      8'b11110111 : _zz_invSub_9 = invSboxRom_247;
      8'b11111000 : _zz_invSub_9 = invSboxRom_248;
      8'b11111001 : _zz_invSub_9 = invSboxRom_249;
      8'b11111010 : _zz_invSub_9 = invSboxRom_250;
      8'b11111011 : _zz_invSub_9 = invSboxRom_251;
      8'b11111100 : _zz_invSub_9 = invSboxRom_252;
      8'b11111101 : _zz_invSub_9 = invSboxRom_253;
      8'b11111110 : _zz_invSub_9 = invSboxRom_254;
      default : _zz_invSub_9 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_10)
      8'b00000000 : _zz_invSub_10 = invSboxRom_0;
      8'b00000001 : _zz_invSub_10 = invSboxRom_1;
      8'b00000010 : _zz_invSub_10 = invSboxRom_2;
      8'b00000011 : _zz_invSub_10 = invSboxRom_3;
      8'b00000100 : _zz_invSub_10 = invSboxRom_4;
      8'b00000101 : _zz_invSub_10 = invSboxRom_5;
      8'b00000110 : _zz_invSub_10 = invSboxRom_6;
      8'b00000111 : _zz_invSub_10 = invSboxRom_7;
      8'b00001000 : _zz_invSub_10 = invSboxRom_8;
      8'b00001001 : _zz_invSub_10 = invSboxRom_9;
      8'b00001010 : _zz_invSub_10 = invSboxRom_10;
      8'b00001011 : _zz_invSub_10 = invSboxRom_11;
      8'b00001100 : _zz_invSub_10 = invSboxRom_12;
      8'b00001101 : _zz_invSub_10 = invSboxRom_13;
      8'b00001110 : _zz_invSub_10 = invSboxRom_14;
      8'b00001111 : _zz_invSub_10 = invSboxRom_15;
      8'b00010000 : _zz_invSub_10 = invSboxRom_16;
      8'b00010001 : _zz_invSub_10 = invSboxRom_17;
      8'b00010010 : _zz_invSub_10 = invSboxRom_18;
      8'b00010011 : _zz_invSub_10 = invSboxRom_19;
      8'b00010100 : _zz_invSub_10 = invSboxRom_20;
      8'b00010101 : _zz_invSub_10 = invSboxRom_21;
      8'b00010110 : _zz_invSub_10 = invSboxRom_22;
      8'b00010111 : _zz_invSub_10 = invSboxRom_23;
      8'b00011000 : _zz_invSub_10 = invSboxRom_24;
      8'b00011001 : _zz_invSub_10 = invSboxRom_25;
      8'b00011010 : _zz_invSub_10 = invSboxRom_26;
      8'b00011011 : _zz_invSub_10 = invSboxRom_27;
      8'b00011100 : _zz_invSub_10 = invSboxRom_28;
      8'b00011101 : _zz_invSub_10 = invSboxRom_29;
      8'b00011110 : _zz_invSub_10 = invSboxRom_30;
      8'b00011111 : _zz_invSub_10 = invSboxRom_31;
      8'b00100000 : _zz_invSub_10 = invSboxRom_32;
      8'b00100001 : _zz_invSub_10 = invSboxRom_33;
      8'b00100010 : _zz_invSub_10 = invSboxRom_34;
      8'b00100011 : _zz_invSub_10 = invSboxRom_35;
      8'b00100100 : _zz_invSub_10 = invSboxRom_36;
      8'b00100101 : _zz_invSub_10 = invSboxRom_37;
      8'b00100110 : _zz_invSub_10 = invSboxRom_38;
      8'b00100111 : _zz_invSub_10 = invSboxRom_39;
      8'b00101000 : _zz_invSub_10 = invSboxRom_40;
      8'b00101001 : _zz_invSub_10 = invSboxRom_41;
      8'b00101010 : _zz_invSub_10 = invSboxRom_42;
      8'b00101011 : _zz_invSub_10 = invSboxRom_43;
      8'b00101100 : _zz_invSub_10 = invSboxRom_44;
      8'b00101101 : _zz_invSub_10 = invSboxRom_45;
      8'b00101110 : _zz_invSub_10 = invSboxRom_46;
      8'b00101111 : _zz_invSub_10 = invSboxRom_47;
      8'b00110000 : _zz_invSub_10 = invSboxRom_48;
      8'b00110001 : _zz_invSub_10 = invSboxRom_49;
      8'b00110010 : _zz_invSub_10 = invSboxRom_50;
      8'b00110011 : _zz_invSub_10 = invSboxRom_51;
      8'b00110100 : _zz_invSub_10 = invSboxRom_52;
      8'b00110101 : _zz_invSub_10 = invSboxRom_53;
      8'b00110110 : _zz_invSub_10 = invSboxRom_54;
      8'b00110111 : _zz_invSub_10 = invSboxRom_55;
      8'b00111000 : _zz_invSub_10 = invSboxRom_56;
      8'b00111001 : _zz_invSub_10 = invSboxRom_57;
      8'b00111010 : _zz_invSub_10 = invSboxRom_58;
      8'b00111011 : _zz_invSub_10 = invSboxRom_59;
      8'b00111100 : _zz_invSub_10 = invSboxRom_60;
      8'b00111101 : _zz_invSub_10 = invSboxRom_61;
      8'b00111110 : _zz_invSub_10 = invSboxRom_62;
      8'b00111111 : _zz_invSub_10 = invSboxRom_63;
      8'b01000000 : _zz_invSub_10 = invSboxRom_64;
      8'b01000001 : _zz_invSub_10 = invSboxRom_65;
      8'b01000010 : _zz_invSub_10 = invSboxRom_66;
      8'b01000011 : _zz_invSub_10 = invSboxRom_67;
      8'b01000100 : _zz_invSub_10 = invSboxRom_68;
      8'b01000101 : _zz_invSub_10 = invSboxRom_69;
      8'b01000110 : _zz_invSub_10 = invSboxRom_70;
      8'b01000111 : _zz_invSub_10 = invSboxRom_71;
      8'b01001000 : _zz_invSub_10 = invSboxRom_72;
      8'b01001001 : _zz_invSub_10 = invSboxRom_73;
      8'b01001010 : _zz_invSub_10 = invSboxRom_74;
      8'b01001011 : _zz_invSub_10 = invSboxRom_75;
      8'b01001100 : _zz_invSub_10 = invSboxRom_76;
      8'b01001101 : _zz_invSub_10 = invSboxRom_77;
      8'b01001110 : _zz_invSub_10 = invSboxRom_78;
      8'b01001111 : _zz_invSub_10 = invSboxRom_79;
      8'b01010000 : _zz_invSub_10 = invSboxRom_80;
      8'b01010001 : _zz_invSub_10 = invSboxRom_81;
      8'b01010010 : _zz_invSub_10 = invSboxRom_82;
      8'b01010011 : _zz_invSub_10 = invSboxRom_83;
      8'b01010100 : _zz_invSub_10 = invSboxRom_84;
      8'b01010101 : _zz_invSub_10 = invSboxRom_85;
      8'b01010110 : _zz_invSub_10 = invSboxRom_86;
      8'b01010111 : _zz_invSub_10 = invSboxRom_87;
      8'b01011000 : _zz_invSub_10 = invSboxRom_88;
      8'b01011001 : _zz_invSub_10 = invSboxRom_89;
      8'b01011010 : _zz_invSub_10 = invSboxRom_90;
      8'b01011011 : _zz_invSub_10 = invSboxRom_91;
      8'b01011100 : _zz_invSub_10 = invSboxRom_92;
      8'b01011101 : _zz_invSub_10 = invSboxRom_93;
      8'b01011110 : _zz_invSub_10 = invSboxRom_94;
      8'b01011111 : _zz_invSub_10 = invSboxRom_95;
      8'b01100000 : _zz_invSub_10 = invSboxRom_96;
      8'b01100001 : _zz_invSub_10 = invSboxRom_97;
      8'b01100010 : _zz_invSub_10 = invSboxRom_98;
      8'b01100011 : _zz_invSub_10 = invSboxRom_99;
      8'b01100100 : _zz_invSub_10 = invSboxRom_100;
      8'b01100101 : _zz_invSub_10 = invSboxRom_101;
      8'b01100110 : _zz_invSub_10 = invSboxRom_102;
      8'b01100111 : _zz_invSub_10 = invSboxRom_103;
      8'b01101000 : _zz_invSub_10 = invSboxRom_104;
      8'b01101001 : _zz_invSub_10 = invSboxRom_105;
      8'b01101010 : _zz_invSub_10 = invSboxRom_106;
      8'b01101011 : _zz_invSub_10 = invSboxRom_107;
      8'b01101100 : _zz_invSub_10 = invSboxRom_108;
      8'b01101101 : _zz_invSub_10 = invSboxRom_109;
      8'b01101110 : _zz_invSub_10 = invSboxRom_110;
      8'b01101111 : _zz_invSub_10 = invSboxRom_111;
      8'b01110000 : _zz_invSub_10 = invSboxRom_112;
      8'b01110001 : _zz_invSub_10 = invSboxRom_113;
      8'b01110010 : _zz_invSub_10 = invSboxRom_114;
      8'b01110011 : _zz_invSub_10 = invSboxRom_115;
      8'b01110100 : _zz_invSub_10 = invSboxRom_116;
      8'b01110101 : _zz_invSub_10 = invSboxRom_117;
      8'b01110110 : _zz_invSub_10 = invSboxRom_118;
      8'b01110111 : _zz_invSub_10 = invSboxRom_119;
      8'b01111000 : _zz_invSub_10 = invSboxRom_120;
      8'b01111001 : _zz_invSub_10 = invSboxRom_121;
      8'b01111010 : _zz_invSub_10 = invSboxRom_122;
      8'b01111011 : _zz_invSub_10 = invSboxRom_123;
      8'b01111100 : _zz_invSub_10 = invSboxRom_124;
      8'b01111101 : _zz_invSub_10 = invSboxRom_125;
      8'b01111110 : _zz_invSub_10 = invSboxRom_126;
      8'b01111111 : _zz_invSub_10 = invSboxRom_127;
      8'b10000000 : _zz_invSub_10 = invSboxRom_128;
      8'b10000001 : _zz_invSub_10 = invSboxRom_129;
      8'b10000010 : _zz_invSub_10 = invSboxRom_130;
      8'b10000011 : _zz_invSub_10 = invSboxRom_131;
      8'b10000100 : _zz_invSub_10 = invSboxRom_132;
      8'b10000101 : _zz_invSub_10 = invSboxRom_133;
      8'b10000110 : _zz_invSub_10 = invSboxRom_134;
      8'b10000111 : _zz_invSub_10 = invSboxRom_135;
      8'b10001000 : _zz_invSub_10 = invSboxRom_136;
      8'b10001001 : _zz_invSub_10 = invSboxRom_137;
      8'b10001010 : _zz_invSub_10 = invSboxRom_138;
      8'b10001011 : _zz_invSub_10 = invSboxRom_139;
      8'b10001100 : _zz_invSub_10 = invSboxRom_140;
      8'b10001101 : _zz_invSub_10 = invSboxRom_141;
      8'b10001110 : _zz_invSub_10 = invSboxRom_142;
      8'b10001111 : _zz_invSub_10 = invSboxRom_143;
      8'b10010000 : _zz_invSub_10 = invSboxRom_144;
      8'b10010001 : _zz_invSub_10 = invSboxRom_145;
      8'b10010010 : _zz_invSub_10 = invSboxRom_146;
      8'b10010011 : _zz_invSub_10 = invSboxRom_147;
      8'b10010100 : _zz_invSub_10 = invSboxRom_148;
      8'b10010101 : _zz_invSub_10 = invSboxRom_149;
      8'b10010110 : _zz_invSub_10 = invSboxRom_150;
      8'b10010111 : _zz_invSub_10 = invSboxRom_151;
      8'b10011000 : _zz_invSub_10 = invSboxRom_152;
      8'b10011001 : _zz_invSub_10 = invSboxRom_153;
      8'b10011010 : _zz_invSub_10 = invSboxRom_154;
      8'b10011011 : _zz_invSub_10 = invSboxRom_155;
      8'b10011100 : _zz_invSub_10 = invSboxRom_156;
      8'b10011101 : _zz_invSub_10 = invSboxRom_157;
      8'b10011110 : _zz_invSub_10 = invSboxRom_158;
      8'b10011111 : _zz_invSub_10 = invSboxRom_159;
      8'b10100000 : _zz_invSub_10 = invSboxRom_160;
      8'b10100001 : _zz_invSub_10 = invSboxRom_161;
      8'b10100010 : _zz_invSub_10 = invSboxRom_162;
      8'b10100011 : _zz_invSub_10 = invSboxRom_163;
      8'b10100100 : _zz_invSub_10 = invSboxRom_164;
      8'b10100101 : _zz_invSub_10 = invSboxRom_165;
      8'b10100110 : _zz_invSub_10 = invSboxRom_166;
      8'b10100111 : _zz_invSub_10 = invSboxRom_167;
      8'b10101000 : _zz_invSub_10 = invSboxRom_168;
      8'b10101001 : _zz_invSub_10 = invSboxRom_169;
      8'b10101010 : _zz_invSub_10 = invSboxRom_170;
      8'b10101011 : _zz_invSub_10 = invSboxRom_171;
      8'b10101100 : _zz_invSub_10 = invSboxRom_172;
      8'b10101101 : _zz_invSub_10 = invSboxRom_173;
      8'b10101110 : _zz_invSub_10 = invSboxRom_174;
      8'b10101111 : _zz_invSub_10 = invSboxRom_175;
      8'b10110000 : _zz_invSub_10 = invSboxRom_176;
      8'b10110001 : _zz_invSub_10 = invSboxRom_177;
      8'b10110010 : _zz_invSub_10 = invSboxRom_178;
      8'b10110011 : _zz_invSub_10 = invSboxRom_179;
      8'b10110100 : _zz_invSub_10 = invSboxRom_180;
      8'b10110101 : _zz_invSub_10 = invSboxRom_181;
      8'b10110110 : _zz_invSub_10 = invSboxRom_182;
      8'b10110111 : _zz_invSub_10 = invSboxRom_183;
      8'b10111000 : _zz_invSub_10 = invSboxRom_184;
      8'b10111001 : _zz_invSub_10 = invSboxRom_185;
      8'b10111010 : _zz_invSub_10 = invSboxRom_186;
      8'b10111011 : _zz_invSub_10 = invSboxRom_187;
      8'b10111100 : _zz_invSub_10 = invSboxRom_188;
      8'b10111101 : _zz_invSub_10 = invSboxRom_189;
      8'b10111110 : _zz_invSub_10 = invSboxRom_190;
      8'b10111111 : _zz_invSub_10 = invSboxRom_191;
      8'b11000000 : _zz_invSub_10 = invSboxRom_192;
      8'b11000001 : _zz_invSub_10 = invSboxRom_193;
      8'b11000010 : _zz_invSub_10 = invSboxRom_194;
      8'b11000011 : _zz_invSub_10 = invSboxRom_195;
      8'b11000100 : _zz_invSub_10 = invSboxRom_196;
      8'b11000101 : _zz_invSub_10 = invSboxRom_197;
      8'b11000110 : _zz_invSub_10 = invSboxRom_198;
      8'b11000111 : _zz_invSub_10 = invSboxRom_199;
      8'b11001000 : _zz_invSub_10 = invSboxRom_200;
      8'b11001001 : _zz_invSub_10 = invSboxRom_201;
      8'b11001010 : _zz_invSub_10 = invSboxRom_202;
      8'b11001011 : _zz_invSub_10 = invSboxRom_203;
      8'b11001100 : _zz_invSub_10 = invSboxRom_204;
      8'b11001101 : _zz_invSub_10 = invSboxRom_205;
      8'b11001110 : _zz_invSub_10 = invSboxRom_206;
      8'b11001111 : _zz_invSub_10 = invSboxRom_207;
      8'b11010000 : _zz_invSub_10 = invSboxRom_208;
      8'b11010001 : _zz_invSub_10 = invSboxRom_209;
      8'b11010010 : _zz_invSub_10 = invSboxRom_210;
      8'b11010011 : _zz_invSub_10 = invSboxRom_211;
      8'b11010100 : _zz_invSub_10 = invSboxRom_212;
      8'b11010101 : _zz_invSub_10 = invSboxRom_213;
      8'b11010110 : _zz_invSub_10 = invSboxRom_214;
      8'b11010111 : _zz_invSub_10 = invSboxRom_215;
      8'b11011000 : _zz_invSub_10 = invSboxRom_216;
      8'b11011001 : _zz_invSub_10 = invSboxRom_217;
      8'b11011010 : _zz_invSub_10 = invSboxRom_218;
      8'b11011011 : _zz_invSub_10 = invSboxRom_219;
      8'b11011100 : _zz_invSub_10 = invSboxRom_220;
      8'b11011101 : _zz_invSub_10 = invSboxRom_221;
      8'b11011110 : _zz_invSub_10 = invSboxRom_222;
      8'b11011111 : _zz_invSub_10 = invSboxRom_223;
      8'b11100000 : _zz_invSub_10 = invSboxRom_224;
      8'b11100001 : _zz_invSub_10 = invSboxRom_225;
      8'b11100010 : _zz_invSub_10 = invSboxRom_226;
      8'b11100011 : _zz_invSub_10 = invSboxRom_227;
      8'b11100100 : _zz_invSub_10 = invSboxRom_228;
      8'b11100101 : _zz_invSub_10 = invSboxRom_229;
      8'b11100110 : _zz_invSub_10 = invSboxRom_230;
      8'b11100111 : _zz_invSub_10 = invSboxRom_231;
      8'b11101000 : _zz_invSub_10 = invSboxRom_232;
      8'b11101001 : _zz_invSub_10 = invSboxRom_233;
      8'b11101010 : _zz_invSub_10 = invSboxRom_234;
      8'b11101011 : _zz_invSub_10 = invSboxRom_235;
      8'b11101100 : _zz_invSub_10 = invSboxRom_236;
      8'b11101101 : _zz_invSub_10 = invSboxRom_237;
      8'b11101110 : _zz_invSub_10 = invSboxRom_238;
      8'b11101111 : _zz_invSub_10 = invSboxRom_239;
      8'b11110000 : _zz_invSub_10 = invSboxRom_240;
      8'b11110001 : _zz_invSub_10 = invSboxRom_241;
      8'b11110010 : _zz_invSub_10 = invSboxRom_242;
      8'b11110011 : _zz_invSub_10 = invSboxRom_243;
      8'b11110100 : _zz_invSub_10 = invSboxRom_244;
      8'b11110101 : _zz_invSub_10 = invSboxRom_245;
      8'b11110110 : _zz_invSub_10 = invSboxRom_246;
      8'b11110111 : _zz_invSub_10 = invSboxRom_247;
      8'b11111000 : _zz_invSub_10 = invSboxRom_248;
      8'b11111001 : _zz_invSub_10 = invSboxRom_249;
      8'b11111010 : _zz_invSub_10 = invSboxRom_250;
      8'b11111011 : _zz_invSub_10 = invSboxRom_251;
      8'b11111100 : _zz_invSub_10 = invSboxRom_252;
      8'b11111101 : _zz_invSub_10 = invSboxRom_253;
      8'b11111110 : _zz_invSub_10 = invSboxRom_254;
      default : _zz_invSub_10 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_11)
      8'b00000000 : _zz_invSub_11 = invSboxRom_0;
      8'b00000001 : _zz_invSub_11 = invSboxRom_1;
      8'b00000010 : _zz_invSub_11 = invSboxRom_2;
      8'b00000011 : _zz_invSub_11 = invSboxRom_3;
      8'b00000100 : _zz_invSub_11 = invSboxRom_4;
      8'b00000101 : _zz_invSub_11 = invSboxRom_5;
      8'b00000110 : _zz_invSub_11 = invSboxRom_6;
      8'b00000111 : _zz_invSub_11 = invSboxRom_7;
      8'b00001000 : _zz_invSub_11 = invSboxRom_8;
      8'b00001001 : _zz_invSub_11 = invSboxRom_9;
      8'b00001010 : _zz_invSub_11 = invSboxRom_10;
      8'b00001011 : _zz_invSub_11 = invSboxRom_11;
      8'b00001100 : _zz_invSub_11 = invSboxRom_12;
      8'b00001101 : _zz_invSub_11 = invSboxRom_13;
      8'b00001110 : _zz_invSub_11 = invSboxRom_14;
      8'b00001111 : _zz_invSub_11 = invSboxRom_15;
      8'b00010000 : _zz_invSub_11 = invSboxRom_16;
      8'b00010001 : _zz_invSub_11 = invSboxRom_17;
      8'b00010010 : _zz_invSub_11 = invSboxRom_18;
      8'b00010011 : _zz_invSub_11 = invSboxRom_19;
      8'b00010100 : _zz_invSub_11 = invSboxRom_20;
      8'b00010101 : _zz_invSub_11 = invSboxRom_21;
      8'b00010110 : _zz_invSub_11 = invSboxRom_22;
      8'b00010111 : _zz_invSub_11 = invSboxRom_23;
      8'b00011000 : _zz_invSub_11 = invSboxRom_24;
      8'b00011001 : _zz_invSub_11 = invSboxRom_25;
      8'b00011010 : _zz_invSub_11 = invSboxRom_26;
      8'b00011011 : _zz_invSub_11 = invSboxRom_27;
      8'b00011100 : _zz_invSub_11 = invSboxRom_28;
      8'b00011101 : _zz_invSub_11 = invSboxRom_29;
      8'b00011110 : _zz_invSub_11 = invSboxRom_30;
      8'b00011111 : _zz_invSub_11 = invSboxRom_31;
      8'b00100000 : _zz_invSub_11 = invSboxRom_32;
      8'b00100001 : _zz_invSub_11 = invSboxRom_33;
      8'b00100010 : _zz_invSub_11 = invSboxRom_34;
      8'b00100011 : _zz_invSub_11 = invSboxRom_35;
      8'b00100100 : _zz_invSub_11 = invSboxRom_36;
      8'b00100101 : _zz_invSub_11 = invSboxRom_37;
      8'b00100110 : _zz_invSub_11 = invSboxRom_38;
      8'b00100111 : _zz_invSub_11 = invSboxRom_39;
      8'b00101000 : _zz_invSub_11 = invSboxRom_40;
      8'b00101001 : _zz_invSub_11 = invSboxRom_41;
      8'b00101010 : _zz_invSub_11 = invSboxRom_42;
      8'b00101011 : _zz_invSub_11 = invSboxRom_43;
      8'b00101100 : _zz_invSub_11 = invSboxRom_44;
      8'b00101101 : _zz_invSub_11 = invSboxRom_45;
      8'b00101110 : _zz_invSub_11 = invSboxRom_46;
      8'b00101111 : _zz_invSub_11 = invSboxRom_47;
      8'b00110000 : _zz_invSub_11 = invSboxRom_48;
      8'b00110001 : _zz_invSub_11 = invSboxRom_49;
      8'b00110010 : _zz_invSub_11 = invSboxRom_50;
      8'b00110011 : _zz_invSub_11 = invSboxRom_51;
      8'b00110100 : _zz_invSub_11 = invSboxRom_52;
      8'b00110101 : _zz_invSub_11 = invSboxRom_53;
      8'b00110110 : _zz_invSub_11 = invSboxRom_54;
      8'b00110111 : _zz_invSub_11 = invSboxRom_55;
      8'b00111000 : _zz_invSub_11 = invSboxRom_56;
      8'b00111001 : _zz_invSub_11 = invSboxRom_57;
      8'b00111010 : _zz_invSub_11 = invSboxRom_58;
      8'b00111011 : _zz_invSub_11 = invSboxRom_59;
      8'b00111100 : _zz_invSub_11 = invSboxRom_60;
      8'b00111101 : _zz_invSub_11 = invSboxRom_61;
      8'b00111110 : _zz_invSub_11 = invSboxRom_62;
      8'b00111111 : _zz_invSub_11 = invSboxRom_63;
      8'b01000000 : _zz_invSub_11 = invSboxRom_64;
      8'b01000001 : _zz_invSub_11 = invSboxRom_65;
      8'b01000010 : _zz_invSub_11 = invSboxRom_66;
      8'b01000011 : _zz_invSub_11 = invSboxRom_67;
      8'b01000100 : _zz_invSub_11 = invSboxRom_68;
      8'b01000101 : _zz_invSub_11 = invSboxRom_69;
      8'b01000110 : _zz_invSub_11 = invSboxRom_70;
      8'b01000111 : _zz_invSub_11 = invSboxRom_71;
      8'b01001000 : _zz_invSub_11 = invSboxRom_72;
      8'b01001001 : _zz_invSub_11 = invSboxRom_73;
      8'b01001010 : _zz_invSub_11 = invSboxRom_74;
      8'b01001011 : _zz_invSub_11 = invSboxRom_75;
      8'b01001100 : _zz_invSub_11 = invSboxRom_76;
      8'b01001101 : _zz_invSub_11 = invSboxRom_77;
      8'b01001110 : _zz_invSub_11 = invSboxRom_78;
      8'b01001111 : _zz_invSub_11 = invSboxRom_79;
      8'b01010000 : _zz_invSub_11 = invSboxRom_80;
      8'b01010001 : _zz_invSub_11 = invSboxRom_81;
      8'b01010010 : _zz_invSub_11 = invSboxRom_82;
      8'b01010011 : _zz_invSub_11 = invSboxRom_83;
      8'b01010100 : _zz_invSub_11 = invSboxRom_84;
      8'b01010101 : _zz_invSub_11 = invSboxRom_85;
      8'b01010110 : _zz_invSub_11 = invSboxRom_86;
      8'b01010111 : _zz_invSub_11 = invSboxRom_87;
      8'b01011000 : _zz_invSub_11 = invSboxRom_88;
      8'b01011001 : _zz_invSub_11 = invSboxRom_89;
      8'b01011010 : _zz_invSub_11 = invSboxRom_90;
      8'b01011011 : _zz_invSub_11 = invSboxRom_91;
      8'b01011100 : _zz_invSub_11 = invSboxRom_92;
      8'b01011101 : _zz_invSub_11 = invSboxRom_93;
      8'b01011110 : _zz_invSub_11 = invSboxRom_94;
      8'b01011111 : _zz_invSub_11 = invSboxRom_95;
      8'b01100000 : _zz_invSub_11 = invSboxRom_96;
      8'b01100001 : _zz_invSub_11 = invSboxRom_97;
      8'b01100010 : _zz_invSub_11 = invSboxRom_98;
      8'b01100011 : _zz_invSub_11 = invSboxRom_99;
      8'b01100100 : _zz_invSub_11 = invSboxRom_100;
      8'b01100101 : _zz_invSub_11 = invSboxRom_101;
      8'b01100110 : _zz_invSub_11 = invSboxRom_102;
      8'b01100111 : _zz_invSub_11 = invSboxRom_103;
      8'b01101000 : _zz_invSub_11 = invSboxRom_104;
      8'b01101001 : _zz_invSub_11 = invSboxRom_105;
      8'b01101010 : _zz_invSub_11 = invSboxRom_106;
      8'b01101011 : _zz_invSub_11 = invSboxRom_107;
      8'b01101100 : _zz_invSub_11 = invSboxRom_108;
      8'b01101101 : _zz_invSub_11 = invSboxRom_109;
      8'b01101110 : _zz_invSub_11 = invSboxRom_110;
      8'b01101111 : _zz_invSub_11 = invSboxRom_111;
      8'b01110000 : _zz_invSub_11 = invSboxRom_112;
      8'b01110001 : _zz_invSub_11 = invSboxRom_113;
      8'b01110010 : _zz_invSub_11 = invSboxRom_114;
      8'b01110011 : _zz_invSub_11 = invSboxRom_115;
      8'b01110100 : _zz_invSub_11 = invSboxRom_116;
      8'b01110101 : _zz_invSub_11 = invSboxRom_117;
      8'b01110110 : _zz_invSub_11 = invSboxRom_118;
      8'b01110111 : _zz_invSub_11 = invSboxRom_119;
      8'b01111000 : _zz_invSub_11 = invSboxRom_120;
      8'b01111001 : _zz_invSub_11 = invSboxRom_121;
      8'b01111010 : _zz_invSub_11 = invSboxRom_122;
      8'b01111011 : _zz_invSub_11 = invSboxRom_123;
      8'b01111100 : _zz_invSub_11 = invSboxRom_124;
      8'b01111101 : _zz_invSub_11 = invSboxRom_125;
      8'b01111110 : _zz_invSub_11 = invSboxRom_126;
      8'b01111111 : _zz_invSub_11 = invSboxRom_127;
      8'b10000000 : _zz_invSub_11 = invSboxRom_128;
      8'b10000001 : _zz_invSub_11 = invSboxRom_129;
      8'b10000010 : _zz_invSub_11 = invSboxRom_130;
      8'b10000011 : _zz_invSub_11 = invSboxRom_131;
      8'b10000100 : _zz_invSub_11 = invSboxRom_132;
      8'b10000101 : _zz_invSub_11 = invSboxRom_133;
      8'b10000110 : _zz_invSub_11 = invSboxRom_134;
      8'b10000111 : _zz_invSub_11 = invSboxRom_135;
      8'b10001000 : _zz_invSub_11 = invSboxRom_136;
      8'b10001001 : _zz_invSub_11 = invSboxRom_137;
      8'b10001010 : _zz_invSub_11 = invSboxRom_138;
      8'b10001011 : _zz_invSub_11 = invSboxRom_139;
      8'b10001100 : _zz_invSub_11 = invSboxRom_140;
      8'b10001101 : _zz_invSub_11 = invSboxRom_141;
      8'b10001110 : _zz_invSub_11 = invSboxRom_142;
      8'b10001111 : _zz_invSub_11 = invSboxRom_143;
      8'b10010000 : _zz_invSub_11 = invSboxRom_144;
      8'b10010001 : _zz_invSub_11 = invSboxRom_145;
      8'b10010010 : _zz_invSub_11 = invSboxRom_146;
      8'b10010011 : _zz_invSub_11 = invSboxRom_147;
      8'b10010100 : _zz_invSub_11 = invSboxRom_148;
      8'b10010101 : _zz_invSub_11 = invSboxRom_149;
      8'b10010110 : _zz_invSub_11 = invSboxRom_150;
      8'b10010111 : _zz_invSub_11 = invSboxRom_151;
      8'b10011000 : _zz_invSub_11 = invSboxRom_152;
      8'b10011001 : _zz_invSub_11 = invSboxRom_153;
      8'b10011010 : _zz_invSub_11 = invSboxRom_154;
      8'b10011011 : _zz_invSub_11 = invSboxRom_155;
      8'b10011100 : _zz_invSub_11 = invSboxRom_156;
      8'b10011101 : _zz_invSub_11 = invSboxRom_157;
      8'b10011110 : _zz_invSub_11 = invSboxRom_158;
      8'b10011111 : _zz_invSub_11 = invSboxRom_159;
      8'b10100000 : _zz_invSub_11 = invSboxRom_160;
      8'b10100001 : _zz_invSub_11 = invSboxRom_161;
      8'b10100010 : _zz_invSub_11 = invSboxRom_162;
      8'b10100011 : _zz_invSub_11 = invSboxRom_163;
      8'b10100100 : _zz_invSub_11 = invSboxRom_164;
      8'b10100101 : _zz_invSub_11 = invSboxRom_165;
      8'b10100110 : _zz_invSub_11 = invSboxRom_166;
      8'b10100111 : _zz_invSub_11 = invSboxRom_167;
      8'b10101000 : _zz_invSub_11 = invSboxRom_168;
      8'b10101001 : _zz_invSub_11 = invSboxRom_169;
      8'b10101010 : _zz_invSub_11 = invSboxRom_170;
      8'b10101011 : _zz_invSub_11 = invSboxRom_171;
      8'b10101100 : _zz_invSub_11 = invSboxRom_172;
      8'b10101101 : _zz_invSub_11 = invSboxRom_173;
      8'b10101110 : _zz_invSub_11 = invSboxRom_174;
      8'b10101111 : _zz_invSub_11 = invSboxRom_175;
      8'b10110000 : _zz_invSub_11 = invSboxRom_176;
      8'b10110001 : _zz_invSub_11 = invSboxRom_177;
      8'b10110010 : _zz_invSub_11 = invSboxRom_178;
      8'b10110011 : _zz_invSub_11 = invSboxRom_179;
      8'b10110100 : _zz_invSub_11 = invSboxRom_180;
      8'b10110101 : _zz_invSub_11 = invSboxRom_181;
      8'b10110110 : _zz_invSub_11 = invSboxRom_182;
      8'b10110111 : _zz_invSub_11 = invSboxRom_183;
      8'b10111000 : _zz_invSub_11 = invSboxRom_184;
      8'b10111001 : _zz_invSub_11 = invSboxRom_185;
      8'b10111010 : _zz_invSub_11 = invSboxRom_186;
      8'b10111011 : _zz_invSub_11 = invSboxRom_187;
      8'b10111100 : _zz_invSub_11 = invSboxRom_188;
      8'b10111101 : _zz_invSub_11 = invSboxRom_189;
      8'b10111110 : _zz_invSub_11 = invSboxRom_190;
      8'b10111111 : _zz_invSub_11 = invSboxRom_191;
      8'b11000000 : _zz_invSub_11 = invSboxRom_192;
      8'b11000001 : _zz_invSub_11 = invSboxRom_193;
      8'b11000010 : _zz_invSub_11 = invSboxRom_194;
      8'b11000011 : _zz_invSub_11 = invSboxRom_195;
      8'b11000100 : _zz_invSub_11 = invSboxRom_196;
      8'b11000101 : _zz_invSub_11 = invSboxRom_197;
      8'b11000110 : _zz_invSub_11 = invSboxRom_198;
      8'b11000111 : _zz_invSub_11 = invSboxRom_199;
      8'b11001000 : _zz_invSub_11 = invSboxRom_200;
      8'b11001001 : _zz_invSub_11 = invSboxRom_201;
      8'b11001010 : _zz_invSub_11 = invSboxRom_202;
      8'b11001011 : _zz_invSub_11 = invSboxRom_203;
      8'b11001100 : _zz_invSub_11 = invSboxRom_204;
      8'b11001101 : _zz_invSub_11 = invSboxRom_205;
      8'b11001110 : _zz_invSub_11 = invSboxRom_206;
      8'b11001111 : _zz_invSub_11 = invSboxRom_207;
      8'b11010000 : _zz_invSub_11 = invSboxRom_208;
      8'b11010001 : _zz_invSub_11 = invSboxRom_209;
      8'b11010010 : _zz_invSub_11 = invSboxRom_210;
      8'b11010011 : _zz_invSub_11 = invSboxRom_211;
      8'b11010100 : _zz_invSub_11 = invSboxRom_212;
      8'b11010101 : _zz_invSub_11 = invSboxRom_213;
      8'b11010110 : _zz_invSub_11 = invSboxRom_214;
      8'b11010111 : _zz_invSub_11 = invSboxRom_215;
      8'b11011000 : _zz_invSub_11 = invSboxRom_216;
      8'b11011001 : _zz_invSub_11 = invSboxRom_217;
      8'b11011010 : _zz_invSub_11 = invSboxRom_218;
      8'b11011011 : _zz_invSub_11 = invSboxRom_219;
      8'b11011100 : _zz_invSub_11 = invSboxRom_220;
      8'b11011101 : _zz_invSub_11 = invSboxRom_221;
      8'b11011110 : _zz_invSub_11 = invSboxRom_222;
      8'b11011111 : _zz_invSub_11 = invSboxRom_223;
      8'b11100000 : _zz_invSub_11 = invSboxRom_224;
      8'b11100001 : _zz_invSub_11 = invSboxRom_225;
      8'b11100010 : _zz_invSub_11 = invSboxRom_226;
      8'b11100011 : _zz_invSub_11 = invSboxRom_227;
      8'b11100100 : _zz_invSub_11 = invSboxRom_228;
      8'b11100101 : _zz_invSub_11 = invSboxRom_229;
      8'b11100110 : _zz_invSub_11 = invSboxRom_230;
      8'b11100111 : _zz_invSub_11 = invSboxRom_231;
      8'b11101000 : _zz_invSub_11 = invSboxRom_232;
      8'b11101001 : _zz_invSub_11 = invSboxRom_233;
      8'b11101010 : _zz_invSub_11 = invSboxRom_234;
      8'b11101011 : _zz_invSub_11 = invSboxRom_235;
      8'b11101100 : _zz_invSub_11 = invSboxRom_236;
      8'b11101101 : _zz_invSub_11 = invSboxRom_237;
      8'b11101110 : _zz_invSub_11 = invSboxRom_238;
      8'b11101111 : _zz_invSub_11 = invSboxRom_239;
      8'b11110000 : _zz_invSub_11 = invSboxRom_240;
      8'b11110001 : _zz_invSub_11 = invSboxRom_241;
      8'b11110010 : _zz_invSub_11 = invSboxRom_242;
      8'b11110011 : _zz_invSub_11 = invSboxRom_243;
      8'b11110100 : _zz_invSub_11 = invSboxRom_244;
      8'b11110101 : _zz_invSub_11 = invSboxRom_245;
      8'b11110110 : _zz_invSub_11 = invSboxRom_246;
      8'b11110111 : _zz_invSub_11 = invSboxRom_247;
      8'b11111000 : _zz_invSub_11 = invSboxRom_248;
      8'b11111001 : _zz_invSub_11 = invSboxRom_249;
      8'b11111010 : _zz_invSub_11 = invSboxRom_250;
      8'b11111011 : _zz_invSub_11 = invSboxRom_251;
      8'b11111100 : _zz_invSub_11 = invSboxRom_252;
      8'b11111101 : _zz_invSub_11 = invSboxRom_253;
      8'b11111110 : _zz_invSub_11 = invSboxRom_254;
      default : _zz_invSub_11 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_12)
      8'b00000000 : _zz_invSub_12 = invSboxRom_0;
      8'b00000001 : _zz_invSub_12 = invSboxRom_1;
      8'b00000010 : _zz_invSub_12 = invSboxRom_2;
      8'b00000011 : _zz_invSub_12 = invSboxRom_3;
      8'b00000100 : _zz_invSub_12 = invSboxRom_4;
      8'b00000101 : _zz_invSub_12 = invSboxRom_5;
      8'b00000110 : _zz_invSub_12 = invSboxRom_6;
      8'b00000111 : _zz_invSub_12 = invSboxRom_7;
      8'b00001000 : _zz_invSub_12 = invSboxRom_8;
      8'b00001001 : _zz_invSub_12 = invSboxRom_9;
      8'b00001010 : _zz_invSub_12 = invSboxRom_10;
      8'b00001011 : _zz_invSub_12 = invSboxRom_11;
      8'b00001100 : _zz_invSub_12 = invSboxRom_12;
      8'b00001101 : _zz_invSub_12 = invSboxRom_13;
      8'b00001110 : _zz_invSub_12 = invSboxRom_14;
      8'b00001111 : _zz_invSub_12 = invSboxRom_15;
      8'b00010000 : _zz_invSub_12 = invSboxRom_16;
      8'b00010001 : _zz_invSub_12 = invSboxRom_17;
      8'b00010010 : _zz_invSub_12 = invSboxRom_18;
      8'b00010011 : _zz_invSub_12 = invSboxRom_19;
      8'b00010100 : _zz_invSub_12 = invSboxRom_20;
      8'b00010101 : _zz_invSub_12 = invSboxRom_21;
      8'b00010110 : _zz_invSub_12 = invSboxRom_22;
      8'b00010111 : _zz_invSub_12 = invSboxRom_23;
      8'b00011000 : _zz_invSub_12 = invSboxRom_24;
      8'b00011001 : _zz_invSub_12 = invSboxRom_25;
      8'b00011010 : _zz_invSub_12 = invSboxRom_26;
      8'b00011011 : _zz_invSub_12 = invSboxRom_27;
      8'b00011100 : _zz_invSub_12 = invSboxRom_28;
      8'b00011101 : _zz_invSub_12 = invSboxRom_29;
      8'b00011110 : _zz_invSub_12 = invSboxRom_30;
      8'b00011111 : _zz_invSub_12 = invSboxRom_31;
      8'b00100000 : _zz_invSub_12 = invSboxRom_32;
      8'b00100001 : _zz_invSub_12 = invSboxRom_33;
      8'b00100010 : _zz_invSub_12 = invSboxRom_34;
      8'b00100011 : _zz_invSub_12 = invSboxRom_35;
      8'b00100100 : _zz_invSub_12 = invSboxRom_36;
      8'b00100101 : _zz_invSub_12 = invSboxRom_37;
      8'b00100110 : _zz_invSub_12 = invSboxRom_38;
      8'b00100111 : _zz_invSub_12 = invSboxRom_39;
      8'b00101000 : _zz_invSub_12 = invSboxRom_40;
      8'b00101001 : _zz_invSub_12 = invSboxRom_41;
      8'b00101010 : _zz_invSub_12 = invSboxRom_42;
      8'b00101011 : _zz_invSub_12 = invSboxRom_43;
      8'b00101100 : _zz_invSub_12 = invSboxRom_44;
      8'b00101101 : _zz_invSub_12 = invSboxRom_45;
      8'b00101110 : _zz_invSub_12 = invSboxRom_46;
      8'b00101111 : _zz_invSub_12 = invSboxRom_47;
      8'b00110000 : _zz_invSub_12 = invSboxRom_48;
      8'b00110001 : _zz_invSub_12 = invSboxRom_49;
      8'b00110010 : _zz_invSub_12 = invSboxRom_50;
      8'b00110011 : _zz_invSub_12 = invSboxRom_51;
      8'b00110100 : _zz_invSub_12 = invSboxRom_52;
      8'b00110101 : _zz_invSub_12 = invSboxRom_53;
      8'b00110110 : _zz_invSub_12 = invSboxRom_54;
      8'b00110111 : _zz_invSub_12 = invSboxRom_55;
      8'b00111000 : _zz_invSub_12 = invSboxRom_56;
      8'b00111001 : _zz_invSub_12 = invSboxRom_57;
      8'b00111010 : _zz_invSub_12 = invSboxRom_58;
      8'b00111011 : _zz_invSub_12 = invSboxRom_59;
      8'b00111100 : _zz_invSub_12 = invSboxRom_60;
      8'b00111101 : _zz_invSub_12 = invSboxRom_61;
      8'b00111110 : _zz_invSub_12 = invSboxRom_62;
      8'b00111111 : _zz_invSub_12 = invSboxRom_63;
      8'b01000000 : _zz_invSub_12 = invSboxRom_64;
      8'b01000001 : _zz_invSub_12 = invSboxRom_65;
      8'b01000010 : _zz_invSub_12 = invSboxRom_66;
      8'b01000011 : _zz_invSub_12 = invSboxRom_67;
      8'b01000100 : _zz_invSub_12 = invSboxRom_68;
      8'b01000101 : _zz_invSub_12 = invSboxRom_69;
      8'b01000110 : _zz_invSub_12 = invSboxRom_70;
      8'b01000111 : _zz_invSub_12 = invSboxRom_71;
      8'b01001000 : _zz_invSub_12 = invSboxRom_72;
      8'b01001001 : _zz_invSub_12 = invSboxRom_73;
      8'b01001010 : _zz_invSub_12 = invSboxRom_74;
      8'b01001011 : _zz_invSub_12 = invSboxRom_75;
      8'b01001100 : _zz_invSub_12 = invSboxRom_76;
      8'b01001101 : _zz_invSub_12 = invSboxRom_77;
      8'b01001110 : _zz_invSub_12 = invSboxRom_78;
      8'b01001111 : _zz_invSub_12 = invSboxRom_79;
      8'b01010000 : _zz_invSub_12 = invSboxRom_80;
      8'b01010001 : _zz_invSub_12 = invSboxRom_81;
      8'b01010010 : _zz_invSub_12 = invSboxRom_82;
      8'b01010011 : _zz_invSub_12 = invSboxRom_83;
      8'b01010100 : _zz_invSub_12 = invSboxRom_84;
      8'b01010101 : _zz_invSub_12 = invSboxRom_85;
      8'b01010110 : _zz_invSub_12 = invSboxRom_86;
      8'b01010111 : _zz_invSub_12 = invSboxRom_87;
      8'b01011000 : _zz_invSub_12 = invSboxRom_88;
      8'b01011001 : _zz_invSub_12 = invSboxRom_89;
      8'b01011010 : _zz_invSub_12 = invSboxRom_90;
      8'b01011011 : _zz_invSub_12 = invSboxRom_91;
      8'b01011100 : _zz_invSub_12 = invSboxRom_92;
      8'b01011101 : _zz_invSub_12 = invSboxRom_93;
      8'b01011110 : _zz_invSub_12 = invSboxRom_94;
      8'b01011111 : _zz_invSub_12 = invSboxRom_95;
      8'b01100000 : _zz_invSub_12 = invSboxRom_96;
      8'b01100001 : _zz_invSub_12 = invSboxRom_97;
      8'b01100010 : _zz_invSub_12 = invSboxRom_98;
      8'b01100011 : _zz_invSub_12 = invSboxRom_99;
      8'b01100100 : _zz_invSub_12 = invSboxRom_100;
      8'b01100101 : _zz_invSub_12 = invSboxRom_101;
      8'b01100110 : _zz_invSub_12 = invSboxRom_102;
      8'b01100111 : _zz_invSub_12 = invSboxRom_103;
      8'b01101000 : _zz_invSub_12 = invSboxRom_104;
      8'b01101001 : _zz_invSub_12 = invSboxRom_105;
      8'b01101010 : _zz_invSub_12 = invSboxRom_106;
      8'b01101011 : _zz_invSub_12 = invSboxRom_107;
      8'b01101100 : _zz_invSub_12 = invSboxRom_108;
      8'b01101101 : _zz_invSub_12 = invSboxRom_109;
      8'b01101110 : _zz_invSub_12 = invSboxRom_110;
      8'b01101111 : _zz_invSub_12 = invSboxRom_111;
      8'b01110000 : _zz_invSub_12 = invSboxRom_112;
      8'b01110001 : _zz_invSub_12 = invSboxRom_113;
      8'b01110010 : _zz_invSub_12 = invSboxRom_114;
      8'b01110011 : _zz_invSub_12 = invSboxRom_115;
      8'b01110100 : _zz_invSub_12 = invSboxRom_116;
      8'b01110101 : _zz_invSub_12 = invSboxRom_117;
      8'b01110110 : _zz_invSub_12 = invSboxRom_118;
      8'b01110111 : _zz_invSub_12 = invSboxRom_119;
      8'b01111000 : _zz_invSub_12 = invSboxRom_120;
      8'b01111001 : _zz_invSub_12 = invSboxRom_121;
      8'b01111010 : _zz_invSub_12 = invSboxRom_122;
      8'b01111011 : _zz_invSub_12 = invSboxRom_123;
      8'b01111100 : _zz_invSub_12 = invSboxRom_124;
      8'b01111101 : _zz_invSub_12 = invSboxRom_125;
      8'b01111110 : _zz_invSub_12 = invSboxRom_126;
      8'b01111111 : _zz_invSub_12 = invSboxRom_127;
      8'b10000000 : _zz_invSub_12 = invSboxRom_128;
      8'b10000001 : _zz_invSub_12 = invSboxRom_129;
      8'b10000010 : _zz_invSub_12 = invSboxRom_130;
      8'b10000011 : _zz_invSub_12 = invSboxRom_131;
      8'b10000100 : _zz_invSub_12 = invSboxRom_132;
      8'b10000101 : _zz_invSub_12 = invSboxRom_133;
      8'b10000110 : _zz_invSub_12 = invSboxRom_134;
      8'b10000111 : _zz_invSub_12 = invSboxRom_135;
      8'b10001000 : _zz_invSub_12 = invSboxRom_136;
      8'b10001001 : _zz_invSub_12 = invSboxRom_137;
      8'b10001010 : _zz_invSub_12 = invSboxRom_138;
      8'b10001011 : _zz_invSub_12 = invSboxRom_139;
      8'b10001100 : _zz_invSub_12 = invSboxRom_140;
      8'b10001101 : _zz_invSub_12 = invSboxRom_141;
      8'b10001110 : _zz_invSub_12 = invSboxRom_142;
      8'b10001111 : _zz_invSub_12 = invSboxRom_143;
      8'b10010000 : _zz_invSub_12 = invSboxRom_144;
      8'b10010001 : _zz_invSub_12 = invSboxRom_145;
      8'b10010010 : _zz_invSub_12 = invSboxRom_146;
      8'b10010011 : _zz_invSub_12 = invSboxRom_147;
      8'b10010100 : _zz_invSub_12 = invSboxRom_148;
      8'b10010101 : _zz_invSub_12 = invSboxRom_149;
      8'b10010110 : _zz_invSub_12 = invSboxRom_150;
      8'b10010111 : _zz_invSub_12 = invSboxRom_151;
      8'b10011000 : _zz_invSub_12 = invSboxRom_152;
      8'b10011001 : _zz_invSub_12 = invSboxRom_153;
      8'b10011010 : _zz_invSub_12 = invSboxRom_154;
      8'b10011011 : _zz_invSub_12 = invSboxRom_155;
      8'b10011100 : _zz_invSub_12 = invSboxRom_156;
      8'b10011101 : _zz_invSub_12 = invSboxRom_157;
      8'b10011110 : _zz_invSub_12 = invSboxRom_158;
      8'b10011111 : _zz_invSub_12 = invSboxRom_159;
      8'b10100000 : _zz_invSub_12 = invSboxRom_160;
      8'b10100001 : _zz_invSub_12 = invSboxRom_161;
      8'b10100010 : _zz_invSub_12 = invSboxRom_162;
      8'b10100011 : _zz_invSub_12 = invSboxRom_163;
      8'b10100100 : _zz_invSub_12 = invSboxRom_164;
      8'b10100101 : _zz_invSub_12 = invSboxRom_165;
      8'b10100110 : _zz_invSub_12 = invSboxRom_166;
      8'b10100111 : _zz_invSub_12 = invSboxRom_167;
      8'b10101000 : _zz_invSub_12 = invSboxRom_168;
      8'b10101001 : _zz_invSub_12 = invSboxRom_169;
      8'b10101010 : _zz_invSub_12 = invSboxRom_170;
      8'b10101011 : _zz_invSub_12 = invSboxRom_171;
      8'b10101100 : _zz_invSub_12 = invSboxRom_172;
      8'b10101101 : _zz_invSub_12 = invSboxRom_173;
      8'b10101110 : _zz_invSub_12 = invSboxRom_174;
      8'b10101111 : _zz_invSub_12 = invSboxRom_175;
      8'b10110000 : _zz_invSub_12 = invSboxRom_176;
      8'b10110001 : _zz_invSub_12 = invSboxRom_177;
      8'b10110010 : _zz_invSub_12 = invSboxRom_178;
      8'b10110011 : _zz_invSub_12 = invSboxRom_179;
      8'b10110100 : _zz_invSub_12 = invSboxRom_180;
      8'b10110101 : _zz_invSub_12 = invSboxRom_181;
      8'b10110110 : _zz_invSub_12 = invSboxRom_182;
      8'b10110111 : _zz_invSub_12 = invSboxRom_183;
      8'b10111000 : _zz_invSub_12 = invSboxRom_184;
      8'b10111001 : _zz_invSub_12 = invSboxRom_185;
      8'b10111010 : _zz_invSub_12 = invSboxRom_186;
      8'b10111011 : _zz_invSub_12 = invSboxRom_187;
      8'b10111100 : _zz_invSub_12 = invSboxRom_188;
      8'b10111101 : _zz_invSub_12 = invSboxRom_189;
      8'b10111110 : _zz_invSub_12 = invSboxRom_190;
      8'b10111111 : _zz_invSub_12 = invSboxRom_191;
      8'b11000000 : _zz_invSub_12 = invSboxRom_192;
      8'b11000001 : _zz_invSub_12 = invSboxRom_193;
      8'b11000010 : _zz_invSub_12 = invSboxRom_194;
      8'b11000011 : _zz_invSub_12 = invSboxRom_195;
      8'b11000100 : _zz_invSub_12 = invSboxRom_196;
      8'b11000101 : _zz_invSub_12 = invSboxRom_197;
      8'b11000110 : _zz_invSub_12 = invSboxRom_198;
      8'b11000111 : _zz_invSub_12 = invSboxRom_199;
      8'b11001000 : _zz_invSub_12 = invSboxRom_200;
      8'b11001001 : _zz_invSub_12 = invSboxRom_201;
      8'b11001010 : _zz_invSub_12 = invSboxRom_202;
      8'b11001011 : _zz_invSub_12 = invSboxRom_203;
      8'b11001100 : _zz_invSub_12 = invSboxRom_204;
      8'b11001101 : _zz_invSub_12 = invSboxRom_205;
      8'b11001110 : _zz_invSub_12 = invSboxRom_206;
      8'b11001111 : _zz_invSub_12 = invSboxRom_207;
      8'b11010000 : _zz_invSub_12 = invSboxRom_208;
      8'b11010001 : _zz_invSub_12 = invSboxRom_209;
      8'b11010010 : _zz_invSub_12 = invSboxRom_210;
      8'b11010011 : _zz_invSub_12 = invSboxRom_211;
      8'b11010100 : _zz_invSub_12 = invSboxRom_212;
      8'b11010101 : _zz_invSub_12 = invSboxRom_213;
      8'b11010110 : _zz_invSub_12 = invSboxRom_214;
      8'b11010111 : _zz_invSub_12 = invSboxRom_215;
      8'b11011000 : _zz_invSub_12 = invSboxRom_216;
      8'b11011001 : _zz_invSub_12 = invSboxRom_217;
      8'b11011010 : _zz_invSub_12 = invSboxRom_218;
      8'b11011011 : _zz_invSub_12 = invSboxRom_219;
      8'b11011100 : _zz_invSub_12 = invSboxRom_220;
      8'b11011101 : _zz_invSub_12 = invSboxRom_221;
      8'b11011110 : _zz_invSub_12 = invSboxRom_222;
      8'b11011111 : _zz_invSub_12 = invSboxRom_223;
      8'b11100000 : _zz_invSub_12 = invSboxRom_224;
      8'b11100001 : _zz_invSub_12 = invSboxRom_225;
      8'b11100010 : _zz_invSub_12 = invSboxRom_226;
      8'b11100011 : _zz_invSub_12 = invSboxRom_227;
      8'b11100100 : _zz_invSub_12 = invSboxRom_228;
      8'b11100101 : _zz_invSub_12 = invSboxRom_229;
      8'b11100110 : _zz_invSub_12 = invSboxRom_230;
      8'b11100111 : _zz_invSub_12 = invSboxRom_231;
      8'b11101000 : _zz_invSub_12 = invSboxRom_232;
      8'b11101001 : _zz_invSub_12 = invSboxRom_233;
      8'b11101010 : _zz_invSub_12 = invSboxRom_234;
      8'b11101011 : _zz_invSub_12 = invSboxRom_235;
      8'b11101100 : _zz_invSub_12 = invSboxRom_236;
      8'b11101101 : _zz_invSub_12 = invSboxRom_237;
      8'b11101110 : _zz_invSub_12 = invSboxRom_238;
      8'b11101111 : _zz_invSub_12 = invSboxRom_239;
      8'b11110000 : _zz_invSub_12 = invSboxRom_240;
      8'b11110001 : _zz_invSub_12 = invSboxRom_241;
      8'b11110010 : _zz_invSub_12 = invSboxRom_242;
      8'b11110011 : _zz_invSub_12 = invSboxRom_243;
      8'b11110100 : _zz_invSub_12 = invSboxRom_244;
      8'b11110101 : _zz_invSub_12 = invSboxRom_245;
      8'b11110110 : _zz_invSub_12 = invSboxRom_246;
      8'b11110111 : _zz_invSub_12 = invSboxRom_247;
      8'b11111000 : _zz_invSub_12 = invSboxRom_248;
      8'b11111001 : _zz_invSub_12 = invSboxRom_249;
      8'b11111010 : _zz_invSub_12 = invSboxRom_250;
      8'b11111011 : _zz_invSub_12 = invSboxRom_251;
      8'b11111100 : _zz_invSub_12 = invSboxRom_252;
      8'b11111101 : _zz_invSub_12 = invSboxRom_253;
      8'b11111110 : _zz_invSub_12 = invSboxRom_254;
      default : _zz_invSub_12 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_13)
      8'b00000000 : _zz_invSub_13 = invSboxRom_0;
      8'b00000001 : _zz_invSub_13 = invSboxRom_1;
      8'b00000010 : _zz_invSub_13 = invSboxRom_2;
      8'b00000011 : _zz_invSub_13 = invSboxRom_3;
      8'b00000100 : _zz_invSub_13 = invSboxRom_4;
      8'b00000101 : _zz_invSub_13 = invSboxRom_5;
      8'b00000110 : _zz_invSub_13 = invSboxRom_6;
      8'b00000111 : _zz_invSub_13 = invSboxRom_7;
      8'b00001000 : _zz_invSub_13 = invSboxRom_8;
      8'b00001001 : _zz_invSub_13 = invSboxRom_9;
      8'b00001010 : _zz_invSub_13 = invSboxRom_10;
      8'b00001011 : _zz_invSub_13 = invSboxRom_11;
      8'b00001100 : _zz_invSub_13 = invSboxRom_12;
      8'b00001101 : _zz_invSub_13 = invSboxRom_13;
      8'b00001110 : _zz_invSub_13 = invSboxRom_14;
      8'b00001111 : _zz_invSub_13 = invSboxRom_15;
      8'b00010000 : _zz_invSub_13 = invSboxRom_16;
      8'b00010001 : _zz_invSub_13 = invSboxRom_17;
      8'b00010010 : _zz_invSub_13 = invSboxRom_18;
      8'b00010011 : _zz_invSub_13 = invSboxRom_19;
      8'b00010100 : _zz_invSub_13 = invSboxRom_20;
      8'b00010101 : _zz_invSub_13 = invSboxRom_21;
      8'b00010110 : _zz_invSub_13 = invSboxRom_22;
      8'b00010111 : _zz_invSub_13 = invSboxRom_23;
      8'b00011000 : _zz_invSub_13 = invSboxRom_24;
      8'b00011001 : _zz_invSub_13 = invSboxRom_25;
      8'b00011010 : _zz_invSub_13 = invSboxRom_26;
      8'b00011011 : _zz_invSub_13 = invSboxRom_27;
      8'b00011100 : _zz_invSub_13 = invSboxRom_28;
      8'b00011101 : _zz_invSub_13 = invSboxRom_29;
      8'b00011110 : _zz_invSub_13 = invSboxRom_30;
      8'b00011111 : _zz_invSub_13 = invSboxRom_31;
      8'b00100000 : _zz_invSub_13 = invSboxRom_32;
      8'b00100001 : _zz_invSub_13 = invSboxRom_33;
      8'b00100010 : _zz_invSub_13 = invSboxRom_34;
      8'b00100011 : _zz_invSub_13 = invSboxRom_35;
      8'b00100100 : _zz_invSub_13 = invSboxRom_36;
      8'b00100101 : _zz_invSub_13 = invSboxRom_37;
      8'b00100110 : _zz_invSub_13 = invSboxRom_38;
      8'b00100111 : _zz_invSub_13 = invSboxRom_39;
      8'b00101000 : _zz_invSub_13 = invSboxRom_40;
      8'b00101001 : _zz_invSub_13 = invSboxRom_41;
      8'b00101010 : _zz_invSub_13 = invSboxRom_42;
      8'b00101011 : _zz_invSub_13 = invSboxRom_43;
      8'b00101100 : _zz_invSub_13 = invSboxRom_44;
      8'b00101101 : _zz_invSub_13 = invSboxRom_45;
      8'b00101110 : _zz_invSub_13 = invSboxRom_46;
      8'b00101111 : _zz_invSub_13 = invSboxRom_47;
      8'b00110000 : _zz_invSub_13 = invSboxRom_48;
      8'b00110001 : _zz_invSub_13 = invSboxRom_49;
      8'b00110010 : _zz_invSub_13 = invSboxRom_50;
      8'b00110011 : _zz_invSub_13 = invSboxRom_51;
      8'b00110100 : _zz_invSub_13 = invSboxRom_52;
      8'b00110101 : _zz_invSub_13 = invSboxRom_53;
      8'b00110110 : _zz_invSub_13 = invSboxRom_54;
      8'b00110111 : _zz_invSub_13 = invSboxRom_55;
      8'b00111000 : _zz_invSub_13 = invSboxRom_56;
      8'b00111001 : _zz_invSub_13 = invSboxRom_57;
      8'b00111010 : _zz_invSub_13 = invSboxRom_58;
      8'b00111011 : _zz_invSub_13 = invSboxRom_59;
      8'b00111100 : _zz_invSub_13 = invSboxRom_60;
      8'b00111101 : _zz_invSub_13 = invSboxRom_61;
      8'b00111110 : _zz_invSub_13 = invSboxRom_62;
      8'b00111111 : _zz_invSub_13 = invSboxRom_63;
      8'b01000000 : _zz_invSub_13 = invSboxRom_64;
      8'b01000001 : _zz_invSub_13 = invSboxRom_65;
      8'b01000010 : _zz_invSub_13 = invSboxRom_66;
      8'b01000011 : _zz_invSub_13 = invSboxRom_67;
      8'b01000100 : _zz_invSub_13 = invSboxRom_68;
      8'b01000101 : _zz_invSub_13 = invSboxRom_69;
      8'b01000110 : _zz_invSub_13 = invSboxRom_70;
      8'b01000111 : _zz_invSub_13 = invSboxRom_71;
      8'b01001000 : _zz_invSub_13 = invSboxRom_72;
      8'b01001001 : _zz_invSub_13 = invSboxRom_73;
      8'b01001010 : _zz_invSub_13 = invSboxRom_74;
      8'b01001011 : _zz_invSub_13 = invSboxRom_75;
      8'b01001100 : _zz_invSub_13 = invSboxRom_76;
      8'b01001101 : _zz_invSub_13 = invSboxRom_77;
      8'b01001110 : _zz_invSub_13 = invSboxRom_78;
      8'b01001111 : _zz_invSub_13 = invSboxRom_79;
      8'b01010000 : _zz_invSub_13 = invSboxRom_80;
      8'b01010001 : _zz_invSub_13 = invSboxRom_81;
      8'b01010010 : _zz_invSub_13 = invSboxRom_82;
      8'b01010011 : _zz_invSub_13 = invSboxRom_83;
      8'b01010100 : _zz_invSub_13 = invSboxRom_84;
      8'b01010101 : _zz_invSub_13 = invSboxRom_85;
      8'b01010110 : _zz_invSub_13 = invSboxRom_86;
      8'b01010111 : _zz_invSub_13 = invSboxRom_87;
      8'b01011000 : _zz_invSub_13 = invSboxRom_88;
      8'b01011001 : _zz_invSub_13 = invSboxRom_89;
      8'b01011010 : _zz_invSub_13 = invSboxRom_90;
      8'b01011011 : _zz_invSub_13 = invSboxRom_91;
      8'b01011100 : _zz_invSub_13 = invSboxRom_92;
      8'b01011101 : _zz_invSub_13 = invSboxRom_93;
      8'b01011110 : _zz_invSub_13 = invSboxRom_94;
      8'b01011111 : _zz_invSub_13 = invSboxRom_95;
      8'b01100000 : _zz_invSub_13 = invSboxRom_96;
      8'b01100001 : _zz_invSub_13 = invSboxRom_97;
      8'b01100010 : _zz_invSub_13 = invSboxRom_98;
      8'b01100011 : _zz_invSub_13 = invSboxRom_99;
      8'b01100100 : _zz_invSub_13 = invSboxRom_100;
      8'b01100101 : _zz_invSub_13 = invSboxRom_101;
      8'b01100110 : _zz_invSub_13 = invSboxRom_102;
      8'b01100111 : _zz_invSub_13 = invSboxRom_103;
      8'b01101000 : _zz_invSub_13 = invSboxRom_104;
      8'b01101001 : _zz_invSub_13 = invSboxRom_105;
      8'b01101010 : _zz_invSub_13 = invSboxRom_106;
      8'b01101011 : _zz_invSub_13 = invSboxRom_107;
      8'b01101100 : _zz_invSub_13 = invSboxRom_108;
      8'b01101101 : _zz_invSub_13 = invSboxRom_109;
      8'b01101110 : _zz_invSub_13 = invSboxRom_110;
      8'b01101111 : _zz_invSub_13 = invSboxRom_111;
      8'b01110000 : _zz_invSub_13 = invSboxRom_112;
      8'b01110001 : _zz_invSub_13 = invSboxRom_113;
      8'b01110010 : _zz_invSub_13 = invSboxRom_114;
      8'b01110011 : _zz_invSub_13 = invSboxRom_115;
      8'b01110100 : _zz_invSub_13 = invSboxRom_116;
      8'b01110101 : _zz_invSub_13 = invSboxRom_117;
      8'b01110110 : _zz_invSub_13 = invSboxRom_118;
      8'b01110111 : _zz_invSub_13 = invSboxRom_119;
      8'b01111000 : _zz_invSub_13 = invSboxRom_120;
      8'b01111001 : _zz_invSub_13 = invSboxRom_121;
      8'b01111010 : _zz_invSub_13 = invSboxRom_122;
      8'b01111011 : _zz_invSub_13 = invSboxRom_123;
      8'b01111100 : _zz_invSub_13 = invSboxRom_124;
      8'b01111101 : _zz_invSub_13 = invSboxRom_125;
      8'b01111110 : _zz_invSub_13 = invSboxRom_126;
      8'b01111111 : _zz_invSub_13 = invSboxRom_127;
      8'b10000000 : _zz_invSub_13 = invSboxRom_128;
      8'b10000001 : _zz_invSub_13 = invSboxRom_129;
      8'b10000010 : _zz_invSub_13 = invSboxRom_130;
      8'b10000011 : _zz_invSub_13 = invSboxRom_131;
      8'b10000100 : _zz_invSub_13 = invSboxRom_132;
      8'b10000101 : _zz_invSub_13 = invSboxRom_133;
      8'b10000110 : _zz_invSub_13 = invSboxRom_134;
      8'b10000111 : _zz_invSub_13 = invSboxRom_135;
      8'b10001000 : _zz_invSub_13 = invSboxRom_136;
      8'b10001001 : _zz_invSub_13 = invSboxRom_137;
      8'b10001010 : _zz_invSub_13 = invSboxRom_138;
      8'b10001011 : _zz_invSub_13 = invSboxRom_139;
      8'b10001100 : _zz_invSub_13 = invSboxRom_140;
      8'b10001101 : _zz_invSub_13 = invSboxRom_141;
      8'b10001110 : _zz_invSub_13 = invSboxRom_142;
      8'b10001111 : _zz_invSub_13 = invSboxRom_143;
      8'b10010000 : _zz_invSub_13 = invSboxRom_144;
      8'b10010001 : _zz_invSub_13 = invSboxRom_145;
      8'b10010010 : _zz_invSub_13 = invSboxRom_146;
      8'b10010011 : _zz_invSub_13 = invSboxRom_147;
      8'b10010100 : _zz_invSub_13 = invSboxRom_148;
      8'b10010101 : _zz_invSub_13 = invSboxRom_149;
      8'b10010110 : _zz_invSub_13 = invSboxRom_150;
      8'b10010111 : _zz_invSub_13 = invSboxRom_151;
      8'b10011000 : _zz_invSub_13 = invSboxRom_152;
      8'b10011001 : _zz_invSub_13 = invSboxRom_153;
      8'b10011010 : _zz_invSub_13 = invSboxRom_154;
      8'b10011011 : _zz_invSub_13 = invSboxRom_155;
      8'b10011100 : _zz_invSub_13 = invSboxRom_156;
      8'b10011101 : _zz_invSub_13 = invSboxRom_157;
      8'b10011110 : _zz_invSub_13 = invSboxRom_158;
      8'b10011111 : _zz_invSub_13 = invSboxRom_159;
      8'b10100000 : _zz_invSub_13 = invSboxRom_160;
      8'b10100001 : _zz_invSub_13 = invSboxRom_161;
      8'b10100010 : _zz_invSub_13 = invSboxRom_162;
      8'b10100011 : _zz_invSub_13 = invSboxRom_163;
      8'b10100100 : _zz_invSub_13 = invSboxRom_164;
      8'b10100101 : _zz_invSub_13 = invSboxRom_165;
      8'b10100110 : _zz_invSub_13 = invSboxRom_166;
      8'b10100111 : _zz_invSub_13 = invSboxRom_167;
      8'b10101000 : _zz_invSub_13 = invSboxRom_168;
      8'b10101001 : _zz_invSub_13 = invSboxRom_169;
      8'b10101010 : _zz_invSub_13 = invSboxRom_170;
      8'b10101011 : _zz_invSub_13 = invSboxRom_171;
      8'b10101100 : _zz_invSub_13 = invSboxRom_172;
      8'b10101101 : _zz_invSub_13 = invSboxRom_173;
      8'b10101110 : _zz_invSub_13 = invSboxRom_174;
      8'b10101111 : _zz_invSub_13 = invSboxRom_175;
      8'b10110000 : _zz_invSub_13 = invSboxRom_176;
      8'b10110001 : _zz_invSub_13 = invSboxRom_177;
      8'b10110010 : _zz_invSub_13 = invSboxRom_178;
      8'b10110011 : _zz_invSub_13 = invSboxRom_179;
      8'b10110100 : _zz_invSub_13 = invSboxRom_180;
      8'b10110101 : _zz_invSub_13 = invSboxRom_181;
      8'b10110110 : _zz_invSub_13 = invSboxRom_182;
      8'b10110111 : _zz_invSub_13 = invSboxRom_183;
      8'b10111000 : _zz_invSub_13 = invSboxRom_184;
      8'b10111001 : _zz_invSub_13 = invSboxRom_185;
      8'b10111010 : _zz_invSub_13 = invSboxRom_186;
      8'b10111011 : _zz_invSub_13 = invSboxRom_187;
      8'b10111100 : _zz_invSub_13 = invSboxRom_188;
      8'b10111101 : _zz_invSub_13 = invSboxRom_189;
      8'b10111110 : _zz_invSub_13 = invSboxRom_190;
      8'b10111111 : _zz_invSub_13 = invSboxRom_191;
      8'b11000000 : _zz_invSub_13 = invSboxRom_192;
      8'b11000001 : _zz_invSub_13 = invSboxRom_193;
      8'b11000010 : _zz_invSub_13 = invSboxRom_194;
      8'b11000011 : _zz_invSub_13 = invSboxRom_195;
      8'b11000100 : _zz_invSub_13 = invSboxRom_196;
      8'b11000101 : _zz_invSub_13 = invSboxRom_197;
      8'b11000110 : _zz_invSub_13 = invSboxRom_198;
      8'b11000111 : _zz_invSub_13 = invSboxRom_199;
      8'b11001000 : _zz_invSub_13 = invSboxRom_200;
      8'b11001001 : _zz_invSub_13 = invSboxRom_201;
      8'b11001010 : _zz_invSub_13 = invSboxRom_202;
      8'b11001011 : _zz_invSub_13 = invSboxRom_203;
      8'b11001100 : _zz_invSub_13 = invSboxRom_204;
      8'b11001101 : _zz_invSub_13 = invSboxRom_205;
      8'b11001110 : _zz_invSub_13 = invSboxRom_206;
      8'b11001111 : _zz_invSub_13 = invSboxRom_207;
      8'b11010000 : _zz_invSub_13 = invSboxRom_208;
      8'b11010001 : _zz_invSub_13 = invSboxRom_209;
      8'b11010010 : _zz_invSub_13 = invSboxRom_210;
      8'b11010011 : _zz_invSub_13 = invSboxRom_211;
      8'b11010100 : _zz_invSub_13 = invSboxRom_212;
      8'b11010101 : _zz_invSub_13 = invSboxRom_213;
      8'b11010110 : _zz_invSub_13 = invSboxRom_214;
      8'b11010111 : _zz_invSub_13 = invSboxRom_215;
      8'b11011000 : _zz_invSub_13 = invSboxRom_216;
      8'b11011001 : _zz_invSub_13 = invSboxRom_217;
      8'b11011010 : _zz_invSub_13 = invSboxRom_218;
      8'b11011011 : _zz_invSub_13 = invSboxRom_219;
      8'b11011100 : _zz_invSub_13 = invSboxRom_220;
      8'b11011101 : _zz_invSub_13 = invSboxRom_221;
      8'b11011110 : _zz_invSub_13 = invSboxRom_222;
      8'b11011111 : _zz_invSub_13 = invSboxRom_223;
      8'b11100000 : _zz_invSub_13 = invSboxRom_224;
      8'b11100001 : _zz_invSub_13 = invSboxRom_225;
      8'b11100010 : _zz_invSub_13 = invSboxRom_226;
      8'b11100011 : _zz_invSub_13 = invSboxRom_227;
      8'b11100100 : _zz_invSub_13 = invSboxRom_228;
      8'b11100101 : _zz_invSub_13 = invSboxRom_229;
      8'b11100110 : _zz_invSub_13 = invSboxRom_230;
      8'b11100111 : _zz_invSub_13 = invSboxRom_231;
      8'b11101000 : _zz_invSub_13 = invSboxRom_232;
      8'b11101001 : _zz_invSub_13 = invSboxRom_233;
      8'b11101010 : _zz_invSub_13 = invSboxRom_234;
      8'b11101011 : _zz_invSub_13 = invSboxRom_235;
      8'b11101100 : _zz_invSub_13 = invSboxRom_236;
      8'b11101101 : _zz_invSub_13 = invSboxRom_237;
      8'b11101110 : _zz_invSub_13 = invSboxRom_238;
      8'b11101111 : _zz_invSub_13 = invSboxRom_239;
      8'b11110000 : _zz_invSub_13 = invSboxRom_240;
      8'b11110001 : _zz_invSub_13 = invSboxRom_241;
      8'b11110010 : _zz_invSub_13 = invSboxRom_242;
      8'b11110011 : _zz_invSub_13 = invSboxRom_243;
      8'b11110100 : _zz_invSub_13 = invSboxRom_244;
      8'b11110101 : _zz_invSub_13 = invSboxRom_245;
      8'b11110110 : _zz_invSub_13 = invSboxRom_246;
      8'b11110111 : _zz_invSub_13 = invSboxRom_247;
      8'b11111000 : _zz_invSub_13 = invSboxRom_248;
      8'b11111001 : _zz_invSub_13 = invSboxRom_249;
      8'b11111010 : _zz_invSub_13 = invSboxRom_250;
      8'b11111011 : _zz_invSub_13 = invSboxRom_251;
      8'b11111100 : _zz_invSub_13 = invSboxRom_252;
      8'b11111101 : _zz_invSub_13 = invSboxRom_253;
      8'b11111110 : _zz_invSub_13 = invSboxRom_254;
      default : _zz_invSub_13 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_14)
      8'b00000000 : _zz_invSub_14 = invSboxRom_0;
      8'b00000001 : _zz_invSub_14 = invSboxRom_1;
      8'b00000010 : _zz_invSub_14 = invSboxRom_2;
      8'b00000011 : _zz_invSub_14 = invSboxRom_3;
      8'b00000100 : _zz_invSub_14 = invSboxRom_4;
      8'b00000101 : _zz_invSub_14 = invSboxRom_5;
      8'b00000110 : _zz_invSub_14 = invSboxRom_6;
      8'b00000111 : _zz_invSub_14 = invSboxRom_7;
      8'b00001000 : _zz_invSub_14 = invSboxRom_8;
      8'b00001001 : _zz_invSub_14 = invSboxRom_9;
      8'b00001010 : _zz_invSub_14 = invSboxRom_10;
      8'b00001011 : _zz_invSub_14 = invSboxRom_11;
      8'b00001100 : _zz_invSub_14 = invSboxRom_12;
      8'b00001101 : _zz_invSub_14 = invSboxRom_13;
      8'b00001110 : _zz_invSub_14 = invSboxRom_14;
      8'b00001111 : _zz_invSub_14 = invSboxRom_15;
      8'b00010000 : _zz_invSub_14 = invSboxRom_16;
      8'b00010001 : _zz_invSub_14 = invSboxRom_17;
      8'b00010010 : _zz_invSub_14 = invSboxRom_18;
      8'b00010011 : _zz_invSub_14 = invSboxRom_19;
      8'b00010100 : _zz_invSub_14 = invSboxRom_20;
      8'b00010101 : _zz_invSub_14 = invSboxRom_21;
      8'b00010110 : _zz_invSub_14 = invSboxRom_22;
      8'b00010111 : _zz_invSub_14 = invSboxRom_23;
      8'b00011000 : _zz_invSub_14 = invSboxRom_24;
      8'b00011001 : _zz_invSub_14 = invSboxRom_25;
      8'b00011010 : _zz_invSub_14 = invSboxRom_26;
      8'b00011011 : _zz_invSub_14 = invSboxRom_27;
      8'b00011100 : _zz_invSub_14 = invSboxRom_28;
      8'b00011101 : _zz_invSub_14 = invSboxRom_29;
      8'b00011110 : _zz_invSub_14 = invSboxRom_30;
      8'b00011111 : _zz_invSub_14 = invSboxRom_31;
      8'b00100000 : _zz_invSub_14 = invSboxRom_32;
      8'b00100001 : _zz_invSub_14 = invSboxRom_33;
      8'b00100010 : _zz_invSub_14 = invSboxRom_34;
      8'b00100011 : _zz_invSub_14 = invSboxRom_35;
      8'b00100100 : _zz_invSub_14 = invSboxRom_36;
      8'b00100101 : _zz_invSub_14 = invSboxRom_37;
      8'b00100110 : _zz_invSub_14 = invSboxRom_38;
      8'b00100111 : _zz_invSub_14 = invSboxRom_39;
      8'b00101000 : _zz_invSub_14 = invSboxRom_40;
      8'b00101001 : _zz_invSub_14 = invSboxRom_41;
      8'b00101010 : _zz_invSub_14 = invSboxRom_42;
      8'b00101011 : _zz_invSub_14 = invSboxRom_43;
      8'b00101100 : _zz_invSub_14 = invSboxRom_44;
      8'b00101101 : _zz_invSub_14 = invSboxRom_45;
      8'b00101110 : _zz_invSub_14 = invSboxRom_46;
      8'b00101111 : _zz_invSub_14 = invSboxRom_47;
      8'b00110000 : _zz_invSub_14 = invSboxRom_48;
      8'b00110001 : _zz_invSub_14 = invSboxRom_49;
      8'b00110010 : _zz_invSub_14 = invSboxRom_50;
      8'b00110011 : _zz_invSub_14 = invSboxRom_51;
      8'b00110100 : _zz_invSub_14 = invSboxRom_52;
      8'b00110101 : _zz_invSub_14 = invSboxRom_53;
      8'b00110110 : _zz_invSub_14 = invSboxRom_54;
      8'b00110111 : _zz_invSub_14 = invSboxRom_55;
      8'b00111000 : _zz_invSub_14 = invSboxRom_56;
      8'b00111001 : _zz_invSub_14 = invSboxRom_57;
      8'b00111010 : _zz_invSub_14 = invSboxRom_58;
      8'b00111011 : _zz_invSub_14 = invSboxRom_59;
      8'b00111100 : _zz_invSub_14 = invSboxRom_60;
      8'b00111101 : _zz_invSub_14 = invSboxRom_61;
      8'b00111110 : _zz_invSub_14 = invSboxRom_62;
      8'b00111111 : _zz_invSub_14 = invSboxRom_63;
      8'b01000000 : _zz_invSub_14 = invSboxRom_64;
      8'b01000001 : _zz_invSub_14 = invSboxRom_65;
      8'b01000010 : _zz_invSub_14 = invSboxRom_66;
      8'b01000011 : _zz_invSub_14 = invSboxRom_67;
      8'b01000100 : _zz_invSub_14 = invSboxRom_68;
      8'b01000101 : _zz_invSub_14 = invSboxRom_69;
      8'b01000110 : _zz_invSub_14 = invSboxRom_70;
      8'b01000111 : _zz_invSub_14 = invSboxRom_71;
      8'b01001000 : _zz_invSub_14 = invSboxRom_72;
      8'b01001001 : _zz_invSub_14 = invSboxRom_73;
      8'b01001010 : _zz_invSub_14 = invSboxRom_74;
      8'b01001011 : _zz_invSub_14 = invSboxRom_75;
      8'b01001100 : _zz_invSub_14 = invSboxRom_76;
      8'b01001101 : _zz_invSub_14 = invSboxRom_77;
      8'b01001110 : _zz_invSub_14 = invSboxRom_78;
      8'b01001111 : _zz_invSub_14 = invSboxRom_79;
      8'b01010000 : _zz_invSub_14 = invSboxRom_80;
      8'b01010001 : _zz_invSub_14 = invSboxRom_81;
      8'b01010010 : _zz_invSub_14 = invSboxRom_82;
      8'b01010011 : _zz_invSub_14 = invSboxRom_83;
      8'b01010100 : _zz_invSub_14 = invSboxRom_84;
      8'b01010101 : _zz_invSub_14 = invSboxRom_85;
      8'b01010110 : _zz_invSub_14 = invSboxRom_86;
      8'b01010111 : _zz_invSub_14 = invSboxRom_87;
      8'b01011000 : _zz_invSub_14 = invSboxRom_88;
      8'b01011001 : _zz_invSub_14 = invSboxRom_89;
      8'b01011010 : _zz_invSub_14 = invSboxRom_90;
      8'b01011011 : _zz_invSub_14 = invSboxRom_91;
      8'b01011100 : _zz_invSub_14 = invSboxRom_92;
      8'b01011101 : _zz_invSub_14 = invSboxRom_93;
      8'b01011110 : _zz_invSub_14 = invSboxRom_94;
      8'b01011111 : _zz_invSub_14 = invSboxRom_95;
      8'b01100000 : _zz_invSub_14 = invSboxRom_96;
      8'b01100001 : _zz_invSub_14 = invSboxRom_97;
      8'b01100010 : _zz_invSub_14 = invSboxRom_98;
      8'b01100011 : _zz_invSub_14 = invSboxRom_99;
      8'b01100100 : _zz_invSub_14 = invSboxRom_100;
      8'b01100101 : _zz_invSub_14 = invSboxRom_101;
      8'b01100110 : _zz_invSub_14 = invSboxRom_102;
      8'b01100111 : _zz_invSub_14 = invSboxRom_103;
      8'b01101000 : _zz_invSub_14 = invSboxRom_104;
      8'b01101001 : _zz_invSub_14 = invSboxRom_105;
      8'b01101010 : _zz_invSub_14 = invSboxRom_106;
      8'b01101011 : _zz_invSub_14 = invSboxRom_107;
      8'b01101100 : _zz_invSub_14 = invSboxRom_108;
      8'b01101101 : _zz_invSub_14 = invSboxRom_109;
      8'b01101110 : _zz_invSub_14 = invSboxRom_110;
      8'b01101111 : _zz_invSub_14 = invSboxRom_111;
      8'b01110000 : _zz_invSub_14 = invSboxRom_112;
      8'b01110001 : _zz_invSub_14 = invSboxRom_113;
      8'b01110010 : _zz_invSub_14 = invSboxRom_114;
      8'b01110011 : _zz_invSub_14 = invSboxRom_115;
      8'b01110100 : _zz_invSub_14 = invSboxRom_116;
      8'b01110101 : _zz_invSub_14 = invSboxRom_117;
      8'b01110110 : _zz_invSub_14 = invSboxRom_118;
      8'b01110111 : _zz_invSub_14 = invSboxRom_119;
      8'b01111000 : _zz_invSub_14 = invSboxRom_120;
      8'b01111001 : _zz_invSub_14 = invSboxRom_121;
      8'b01111010 : _zz_invSub_14 = invSboxRom_122;
      8'b01111011 : _zz_invSub_14 = invSboxRom_123;
      8'b01111100 : _zz_invSub_14 = invSboxRom_124;
      8'b01111101 : _zz_invSub_14 = invSboxRom_125;
      8'b01111110 : _zz_invSub_14 = invSboxRom_126;
      8'b01111111 : _zz_invSub_14 = invSboxRom_127;
      8'b10000000 : _zz_invSub_14 = invSboxRom_128;
      8'b10000001 : _zz_invSub_14 = invSboxRom_129;
      8'b10000010 : _zz_invSub_14 = invSboxRom_130;
      8'b10000011 : _zz_invSub_14 = invSboxRom_131;
      8'b10000100 : _zz_invSub_14 = invSboxRom_132;
      8'b10000101 : _zz_invSub_14 = invSboxRom_133;
      8'b10000110 : _zz_invSub_14 = invSboxRom_134;
      8'b10000111 : _zz_invSub_14 = invSboxRom_135;
      8'b10001000 : _zz_invSub_14 = invSboxRom_136;
      8'b10001001 : _zz_invSub_14 = invSboxRom_137;
      8'b10001010 : _zz_invSub_14 = invSboxRom_138;
      8'b10001011 : _zz_invSub_14 = invSboxRom_139;
      8'b10001100 : _zz_invSub_14 = invSboxRom_140;
      8'b10001101 : _zz_invSub_14 = invSboxRom_141;
      8'b10001110 : _zz_invSub_14 = invSboxRom_142;
      8'b10001111 : _zz_invSub_14 = invSboxRom_143;
      8'b10010000 : _zz_invSub_14 = invSboxRom_144;
      8'b10010001 : _zz_invSub_14 = invSboxRom_145;
      8'b10010010 : _zz_invSub_14 = invSboxRom_146;
      8'b10010011 : _zz_invSub_14 = invSboxRom_147;
      8'b10010100 : _zz_invSub_14 = invSboxRom_148;
      8'b10010101 : _zz_invSub_14 = invSboxRom_149;
      8'b10010110 : _zz_invSub_14 = invSboxRom_150;
      8'b10010111 : _zz_invSub_14 = invSboxRom_151;
      8'b10011000 : _zz_invSub_14 = invSboxRom_152;
      8'b10011001 : _zz_invSub_14 = invSboxRom_153;
      8'b10011010 : _zz_invSub_14 = invSboxRom_154;
      8'b10011011 : _zz_invSub_14 = invSboxRom_155;
      8'b10011100 : _zz_invSub_14 = invSboxRom_156;
      8'b10011101 : _zz_invSub_14 = invSboxRom_157;
      8'b10011110 : _zz_invSub_14 = invSboxRom_158;
      8'b10011111 : _zz_invSub_14 = invSboxRom_159;
      8'b10100000 : _zz_invSub_14 = invSboxRom_160;
      8'b10100001 : _zz_invSub_14 = invSboxRom_161;
      8'b10100010 : _zz_invSub_14 = invSboxRom_162;
      8'b10100011 : _zz_invSub_14 = invSboxRom_163;
      8'b10100100 : _zz_invSub_14 = invSboxRom_164;
      8'b10100101 : _zz_invSub_14 = invSboxRom_165;
      8'b10100110 : _zz_invSub_14 = invSboxRom_166;
      8'b10100111 : _zz_invSub_14 = invSboxRom_167;
      8'b10101000 : _zz_invSub_14 = invSboxRom_168;
      8'b10101001 : _zz_invSub_14 = invSboxRom_169;
      8'b10101010 : _zz_invSub_14 = invSboxRom_170;
      8'b10101011 : _zz_invSub_14 = invSboxRom_171;
      8'b10101100 : _zz_invSub_14 = invSboxRom_172;
      8'b10101101 : _zz_invSub_14 = invSboxRom_173;
      8'b10101110 : _zz_invSub_14 = invSboxRom_174;
      8'b10101111 : _zz_invSub_14 = invSboxRom_175;
      8'b10110000 : _zz_invSub_14 = invSboxRom_176;
      8'b10110001 : _zz_invSub_14 = invSboxRom_177;
      8'b10110010 : _zz_invSub_14 = invSboxRom_178;
      8'b10110011 : _zz_invSub_14 = invSboxRom_179;
      8'b10110100 : _zz_invSub_14 = invSboxRom_180;
      8'b10110101 : _zz_invSub_14 = invSboxRom_181;
      8'b10110110 : _zz_invSub_14 = invSboxRom_182;
      8'b10110111 : _zz_invSub_14 = invSboxRom_183;
      8'b10111000 : _zz_invSub_14 = invSboxRom_184;
      8'b10111001 : _zz_invSub_14 = invSboxRom_185;
      8'b10111010 : _zz_invSub_14 = invSboxRom_186;
      8'b10111011 : _zz_invSub_14 = invSboxRom_187;
      8'b10111100 : _zz_invSub_14 = invSboxRom_188;
      8'b10111101 : _zz_invSub_14 = invSboxRom_189;
      8'b10111110 : _zz_invSub_14 = invSboxRom_190;
      8'b10111111 : _zz_invSub_14 = invSboxRom_191;
      8'b11000000 : _zz_invSub_14 = invSboxRom_192;
      8'b11000001 : _zz_invSub_14 = invSboxRom_193;
      8'b11000010 : _zz_invSub_14 = invSboxRom_194;
      8'b11000011 : _zz_invSub_14 = invSboxRom_195;
      8'b11000100 : _zz_invSub_14 = invSboxRom_196;
      8'b11000101 : _zz_invSub_14 = invSboxRom_197;
      8'b11000110 : _zz_invSub_14 = invSboxRom_198;
      8'b11000111 : _zz_invSub_14 = invSboxRom_199;
      8'b11001000 : _zz_invSub_14 = invSboxRom_200;
      8'b11001001 : _zz_invSub_14 = invSboxRom_201;
      8'b11001010 : _zz_invSub_14 = invSboxRom_202;
      8'b11001011 : _zz_invSub_14 = invSboxRom_203;
      8'b11001100 : _zz_invSub_14 = invSboxRom_204;
      8'b11001101 : _zz_invSub_14 = invSboxRom_205;
      8'b11001110 : _zz_invSub_14 = invSboxRom_206;
      8'b11001111 : _zz_invSub_14 = invSboxRom_207;
      8'b11010000 : _zz_invSub_14 = invSboxRom_208;
      8'b11010001 : _zz_invSub_14 = invSboxRom_209;
      8'b11010010 : _zz_invSub_14 = invSboxRom_210;
      8'b11010011 : _zz_invSub_14 = invSboxRom_211;
      8'b11010100 : _zz_invSub_14 = invSboxRom_212;
      8'b11010101 : _zz_invSub_14 = invSboxRom_213;
      8'b11010110 : _zz_invSub_14 = invSboxRom_214;
      8'b11010111 : _zz_invSub_14 = invSboxRom_215;
      8'b11011000 : _zz_invSub_14 = invSboxRom_216;
      8'b11011001 : _zz_invSub_14 = invSboxRom_217;
      8'b11011010 : _zz_invSub_14 = invSboxRom_218;
      8'b11011011 : _zz_invSub_14 = invSboxRom_219;
      8'b11011100 : _zz_invSub_14 = invSboxRom_220;
      8'b11011101 : _zz_invSub_14 = invSboxRom_221;
      8'b11011110 : _zz_invSub_14 = invSboxRom_222;
      8'b11011111 : _zz_invSub_14 = invSboxRom_223;
      8'b11100000 : _zz_invSub_14 = invSboxRom_224;
      8'b11100001 : _zz_invSub_14 = invSboxRom_225;
      8'b11100010 : _zz_invSub_14 = invSboxRom_226;
      8'b11100011 : _zz_invSub_14 = invSboxRom_227;
      8'b11100100 : _zz_invSub_14 = invSboxRom_228;
      8'b11100101 : _zz_invSub_14 = invSboxRom_229;
      8'b11100110 : _zz_invSub_14 = invSboxRom_230;
      8'b11100111 : _zz_invSub_14 = invSboxRom_231;
      8'b11101000 : _zz_invSub_14 = invSboxRom_232;
      8'b11101001 : _zz_invSub_14 = invSboxRom_233;
      8'b11101010 : _zz_invSub_14 = invSboxRom_234;
      8'b11101011 : _zz_invSub_14 = invSboxRom_235;
      8'b11101100 : _zz_invSub_14 = invSboxRom_236;
      8'b11101101 : _zz_invSub_14 = invSboxRom_237;
      8'b11101110 : _zz_invSub_14 = invSboxRom_238;
      8'b11101111 : _zz_invSub_14 = invSboxRom_239;
      8'b11110000 : _zz_invSub_14 = invSboxRom_240;
      8'b11110001 : _zz_invSub_14 = invSboxRom_241;
      8'b11110010 : _zz_invSub_14 = invSboxRom_242;
      8'b11110011 : _zz_invSub_14 = invSboxRom_243;
      8'b11110100 : _zz_invSub_14 = invSboxRom_244;
      8'b11110101 : _zz_invSub_14 = invSboxRom_245;
      8'b11110110 : _zz_invSub_14 = invSboxRom_246;
      8'b11110111 : _zz_invSub_14 = invSboxRom_247;
      8'b11111000 : _zz_invSub_14 = invSboxRom_248;
      8'b11111001 : _zz_invSub_14 = invSboxRom_249;
      8'b11111010 : _zz_invSub_14 = invSboxRom_250;
      8'b11111011 : _zz_invSub_14 = invSboxRom_251;
      8'b11111100 : _zz_invSub_14 = invSboxRom_252;
      8'b11111101 : _zz_invSub_14 = invSboxRom_253;
      8'b11111110 : _zz_invSub_14 = invSboxRom_254;
      default : _zz_invSub_14 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(invShifted_15)
      8'b00000000 : _zz_invSub_15 = invSboxRom_0;
      8'b00000001 : _zz_invSub_15 = invSboxRom_1;
      8'b00000010 : _zz_invSub_15 = invSboxRom_2;
      8'b00000011 : _zz_invSub_15 = invSboxRom_3;
      8'b00000100 : _zz_invSub_15 = invSboxRom_4;
      8'b00000101 : _zz_invSub_15 = invSboxRom_5;
      8'b00000110 : _zz_invSub_15 = invSboxRom_6;
      8'b00000111 : _zz_invSub_15 = invSboxRom_7;
      8'b00001000 : _zz_invSub_15 = invSboxRom_8;
      8'b00001001 : _zz_invSub_15 = invSboxRom_9;
      8'b00001010 : _zz_invSub_15 = invSboxRom_10;
      8'b00001011 : _zz_invSub_15 = invSboxRom_11;
      8'b00001100 : _zz_invSub_15 = invSboxRom_12;
      8'b00001101 : _zz_invSub_15 = invSboxRom_13;
      8'b00001110 : _zz_invSub_15 = invSboxRom_14;
      8'b00001111 : _zz_invSub_15 = invSboxRom_15;
      8'b00010000 : _zz_invSub_15 = invSboxRom_16;
      8'b00010001 : _zz_invSub_15 = invSboxRom_17;
      8'b00010010 : _zz_invSub_15 = invSboxRom_18;
      8'b00010011 : _zz_invSub_15 = invSboxRom_19;
      8'b00010100 : _zz_invSub_15 = invSboxRom_20;
      8'b00010101 : _zz_invSub_15 = invSboxRom_21;
      8'b00010110 : _zz_invSub_15 = invSboxRom_22;
      8'b00010111 : _zz_invSub_15 = invSboxRom_23;
      8'b00011000 : _zz_invSub_15 = invSboxRom_24;
      8'b00011001 : _zz_invSub_15 = invSboxRom_25;
      8'b00011010 : _zz_invSub_15 = invSboxRom_26;
      8'b00011011 : _zz_invSub_15 = invSboxRom_27;
      8'b00011100 : _zz_invSub_15 = invSboxRom_28;
      8'b00011101 : _zz_invSub_15 = invSboxRom_29;
      8'b00011110 : _zz_invSub_15 = invSboxRom_30;
      8'b00011111 : _zz_invSub_15 = invSboxRom_31;
      8'b00100000 : _zz_invSub_15 = invSboxRom_32;
      8'b00100001 : _zz_invSub_15 = invSboxRom_33;
      8'b00100010 : _zz_invSub_15 = invSboxRom_34;
      8'b00100011 : _zz_invSub_15 = invSboxRom_35;
      8'b00100100 : _zz_invSub_15 = invSboxRom_36;
      8'b00100101 : _zz_invSub_15 = invSboxRom_37;
      8'b00100110 : _zz_invSub_15 = invSboxRom_38;
      8'b00100111 : _zz_invSub_15 = invSboxRom_39;
      8'b00101000 : _zz_invSub_15 = invSboxRom_40;
      8'b00101001 : _zz_invSub_15 = invSboxRom_41;
      8'b00101010 : _zz_invSub_15 = invSboxRom_42;
      8'b00101011 : _zz_invSub_15 = invSboxRom_43;
      8'b00101100 : _zz_invSub_15 = invSboxRom_44;
      8'b00101101 : _zz_invSub_15 = invSboxRom_45;
      8'b00101110 : _zz_invSub_15 = invSboxRom_46;
      8'b00101111 : _zz_invSub_15 = invSboxRom_47;
      8'b00110000 : _zz_invSub_15 = invSboxRom_48;
      8'b00110001 : _zz_invSub_15 = invSboxRom_49;
      8'b00110010 : _zz_invSub_15 = invSboxRom_50;
      8'b00110011 : _zz_invSub_15 = invSboxRom_51;
      8'b00110100 : _zz_invSub_15 = invSboxRom_52;
      8'b00110101 : _zz_invSub_15 = invSboxRom_53;
      8'b00110110 : _zz_invSub_15 = invSboxRom_54;
      8'b00110111 : _zz_invSub_15 = invSboxRom_55;
      8'b00111000 : _zz_invSub_15 = invSboxRom_56;
      8'b00111001 : _zz_invSub_15 = invSboxRom_57;
      8'b00111010 : _zz_invSub_15 = invSboxRom_58;
      8'b00111011 : _zz_invSub_15 = invSboxRom_59;
      8'b00111100 : _zz_invSub_15 = invSboxRom_60;
      8'b00111101 : _zz_invSub_15 = invSboxRom_61;
      8'b00111110 : _zz_invSub_15 = invSboxRom_62;
      8'b00111111 : _zz_invSub_15 = invSboxRom_63;
      8'b01000000 : _zz_invSub_15 = invSboxRom_64;
      8'b01000001 : _zz_invSub_15 = invSboxRom_65;
      8'b01000010 : _zz_invSub_15 = invSboxRom_66;
      8'b01000011 : _zz_invSub_15 = invSboxRom_67;
      8'b01000100 : _zz_invSub_15 = invSboxRom_68;
      8'b01000101 : _zz_invSub_15 = invSboxRom_69;
      8'b01000110 : _zz_invSub_15 = invSboxRom_70;
      8'b01000111 : _zz_invSub_15 = invSboxRom_71;
      8'b01001000 : _zz_invSub_15 = invSboxRom_72;
      8'b01001001 : _zz_invSub_15 = invSboxRom_73;
      8'b01001010 : _zz_invSub_15 = invSboxRom_74;
      8'b01001011 : _zz_invSub_15 = invSboxRom_75;
      8'b01001100 : _zz_invSub_15 = invSboxRom_76;
      8'b01001101 : _zz_invSub_15 = invSboxRom_77;
      8'b01001110 : _zz_invSub_15 = invSboxRom_78;
      8'b01001111 : _zz_invSub_15 = invSboxRom_79;
      8'b01010000 : _zz_invSub_15 = invSboxRom_80;
      8'b01010001 : _zz_invSub_15 = invSboxRom_81;
      8'b01010010 : _zz_invSub_15 = invSboxRom_82;
      8'b01010011 : _zz_invSub_15 = invSboxRom_83;
      8'b01010100 : _zz_invSub_15 = invSboxRom_84;
      8'b01010101 : _zz_invSub_15 = invSboxRom_85;
      8'b01010110 : _zz_invSub_15 = invSboxRom_86;
      8'b01010111 : _zz_invSub_15 = invSboxRom_87;
      8'b01011000 : _zz_invSub_15 = invSboxRom_88;
      8'b01011001 : _zz_invSub_15 = invSboxRom_89;
      8'b01011010 : _zz_invSub_15 = invSboxRom_90;
      8'b01011011 : _zz_invSub_15 = invSboxRom_91;
      8'b01011100 : _zz_invSub_15 = invSboxRom_92;
      8'b01011101 : _zz_invSub_15 = invSboxRom_93;
      8'b01011110 : _zz_invSub_15 = invSboxRom_94;
      8'b01011111 : _zz_invSub_15 = invSboxRom_95;
      8'b01100000 : _zz_invSub_15 = invSboxRom_96;
      8'b01100001 : _zz_invSub_15 = invSboxRom_97;
      8'b01100010 : _zz_invSub_15 = invSboxRom_98;
      8'b01100011 : _zz_invSub_15 = invSboxRom_99;
      8'b01100100 : _zz_invSub_15 = invSboxRom_100;
      8'b01100101 : _zz_invSub_15 = invSboxRom_101;
      8'b01100110 : _zz_invSub_15 = invSboxRom_102;
      8'b01100111 : _zz_invSub_15 = invSboxRom_103;
      8'b01101000 : _zz_invSub_15 = invSboxRom_104;
      8'b01101001 : _zz_invSub_15 = invSboxRom_105;
      8'b01101010 : _zz_invSub_15 = invSboxRom_106;
      8'b01101011 : _zz_invSub_15 = invSboxRom_107;
      8'b01101100 : _zz_invSub_15 = invSboxRom_108;
      8'b01101101 : _zz_invSub_15 = invSboxRom_109;
      8'b01101110 : _zz_invSub_15 = invSboxRom_110;
      8'b01101111 : _zz_invSub_15 = invSboxRom_111;
      8'b01110000 : _zz_invSub_15 = invSboxRom_112;
      8'b01110001 : _zz_invSub_15 = invSboxRom_113;
      8'b01110010 : _zz_invSub_15 = invSboxRom_114;
      8'b01110011 : _zz_invSub_15 = invSboxRom_115;
      8'b01110100 : _zz_invSub_15 = invSboxRom_116;
      8'b01110101 : _zz_invSub_15 = invSboxRom_117;
      8'b01110110 : _zz_invSub_15 = invSboxRom_118;
      8'b01110111 : _zz_invSub_15 = invSboxRom_119;
      8'b01111000 : _zz_invSub_15 = invSboxRom_120;
      8'b01111001 : _zz_invSub_15 = invSboxRom_121;
      8'b01111010 : _zz_invSub_15 = invSboxRom_122;
      8'b01111011 : _zz_invSub_15 = invSboxRom_123;
      8'b01111100 : _zz_invSub_15 = invSboxRom_124;
      8'b01111101 : _zz_invSub_15 = invSboxRom_125;
      8'b01111110 : _zz_invSub_15 = invSboxRom_126;
      8'b01111111 : _zz_invSub_15 = invSboxRom_127;
      8'b10000000 : _zz_invSub_15 = invSboxRom_128;
      8'b10000001 : _zz_invSub_15 = invSboxRom_129;
      8'b10000010 : _zz_invSub_15 = invSboxRom_130;
      8'b10000011 : _zz_invSub_15 = invSboxRom_131;
      8'b10000100 : _zz_invSub_15 = invSboxRom_132;
      8'b10000101 : _zz_invSub_15 = invSboxRom_133;
      8'b10000110 : _zz_invSub_15 = invSboxRom_134;
      8'b10000111 : _zz_invSub_15 = invSboxRom_135;
      8'b10001000 : _zz_invSub_15 = invSboxRom_136;
      8'b10001001 : _zz_invSub_15 = invSboxRom_137;
      8'b10001010 : _zz_invSub_15 = invSboxRom_138;
      8'b10001011 : _zz_invSub_15 = invSboxRom_139;
      8'b10001100 : _zz_invSub_15 = invSboxRom_140;
      8'b10001101 : _zz_invSub_15 = invSboxRom_141;
      8'b10001110 : _zz_invSub_15 = invSboxRom_142;
      8'b10001111 : _zz_invSub_15 = invSboxRom_143;
      8'b10010000 : _zz_invSub_15 = invSboxRom_144;
      8'b10010001 : _zz_invSub_15 = invSboxRom_145;
      8'b10010010 : _zz_invSub_15 = invSboxRom_146;
      8'b10010011 : _zz_invSub_15 = invSboxRom_147;
      8'b10010100 : _zz_invSub_15 = invSboxRom_148;
      8'b10010101 : _zz_invSub_15 = invSboxRom_149;
      8'b10010110 : _zz_invSub_15 = invSboxRom_150;
      8'b10010111 : _zz_invSub_15 = invSboxRom_151;
      8'b10011000 : _zz_invSub_15 = invSboxRom_152;
      8'b10011001 : _zz_invSub_15 = invSboxRom_153;
      8'b10011010 : _zz_invSub_15 = invSboxRom_154;
      8'b10011011 : _zz_invSub_15 = invSboxRom_155;
      8'b10011100 : _zz_invSub_15 = invSboxRom_156;
      8'b10011101 : _zz_invSub_15 = invSboxRom_157;
      8'b10011110 : _zz_invSub_15 = invSboxRom_158;
      8'b10011111 : _zz_invSub_15 = invSboxRom_159;
      8'b10100000 : _zz_invSub_15 = invSboxRom_160;
      8'b10100001 : _zz_invSub_15 = invSboxRom_161;
      8'b10100010 : _zz_invSub_15 = invSboxRom_162;
      8'b10100011 : _zz_invSub_15 = invSboxRom_163;
      8'b10100100 : _zz_invSub_15 = invSboxRom_164;
      8'b10100101 : _zz_invSub_15 = invSboxRom_165;
      8'b10100110 : _zz_invSub_15 = invSboxRom_166;
      8'b10100111 : _zz_invSub_15 = invSboxRom_167;
      8'b10101000 : _zz_invSub_15 = invSboxRom_168;
      8'b10101001 : _zz_invSub_15 = invSboxRom_169;
      8'b10101010 : _zz_invSub_15 = invSboxRom_170;
      8'b10101011 : _zz_invSub_15 = invSboxRom_171;
      8'b10101100 : _zz_invSub_15 = invSboxRom_172;
      8'b10101101 : _zz_invSub_15 = invSboxRom_173;
      8'b10101110 : _zz_invSub_15 = invSboxRom_174;
      8'b10101111 : _zz_invSub_15 = invSboxRom_175;
      8'b10110000 : _zz_invSub_15 = invSboxRom_176;
      8'b10110001 : _zz_invSub_15 = invSboxRom_177;
      8'b10110010 : _zz_invSub_15 = invSboxRom_178;
      8'b10110011 : _zz_invSub_15 = invSboxRom_179;
      8'b10110100 : _zz_invSub_15 = invSboxRom_180;
      8'b10110101 : _zz_invSub_15 = invSboxRom_181;
      8'b10110110 : _zz_invSub_15 = invSboxRom_182;
      8'b10110111 : _zz_invSub_15 = invSboxRom_183;
      8'b10111000 : _zz_invSub_15 = invSboxRom_184;
      8'b10111001 : _zz_invSub_15 = invSboxRom_185;
      8'b10111010 : _zz_invSub_15 = invSboxRom_186;
      8'b10111011 : _zz_invSub_15 = invSboxRom_187;
      8'b10111100 : _zz_invSub_15 = invSboxRom_188;
      8'b10111101 : _zz_invSub_15 = invSboxRom_189;
      8'b10111110 : _zz_invSub_15 = invSboxRom_190;
      8'b10111111 : _zz_invSub_15 = invSboxRom_191;
      8'b11000000 : _zz_invSub_15 = invSboxRom_192;
      8'b11000001 : _zz_invSub_15 = invSboxRom_193;
      8'b11000010 : _zz_invSub_15 = invSboxRom_194;
      8'b11000011 : _zz_invSub_15 = invSboxRom_195;
      8'b11000100 : _zz_invSub_15 = invSboxRom_196;
      8'b11000101 : _zz_invSub_15 = invSboxRom_197;
      8'b11000110 : _zz_invSub_15 = invSboxRom_198;
      8'b11000111 : _zz_invSub_15 = invSboxRom_199;
      8'b11001000 : _zz_invSub_15 = invSboxRom_200;
      8'b11001001 : _zz_invSub_15 = invSboxRom_201;
      8'b11001010 : _zz_invSub_15 = invSboxRom_202;
      8'b11001011 : _zz_invSub_15 = invSboxRom_203;
      8'b11001100 : _zz_invSub_15 = invSboxRom_204;
      8'b11001101 : _zz_invSub_15 = invSboxRom_205;
      8'b11001110 : _zz_invSub_15 = invSboxRom_206;
      8'b11001111 : _zz_invSub_15 = invSboxRom_207;
      8'b11010000 : _zz_invSub_15 = invSboxRom_208;
      8'b11010001 : _zz_invSub_15 = invSboxRom_209;
      8'b11010010 : _zz_invSub_15 = invSboxRom_210;
      8'b11010011 : _zz_invSub_15 = invSboxRom_211;
      8'b11010100 : _zz_invSub_15 = invSboxRom_212;
      8'b11010101 : _zz_invSub_15 = invSboxRom_213;
      8'b11010110 : _zz_invSub_15 = invSboxRom_214;
      8'b11010111 : _zz_invSub_15 = invSboxRom_215;
      8'b11011000 : _zz_invSub_15 = invSboxRom_216;
      8'b11011001 : _zz_invSub_15 = invSboxRom_217;
      8'b11011010 : _zz_invSub_15 = invSboxRom_218;
      8'b11011011 : _zz_invSub_15 = invSboxRom_219;
      8'b11011100 : _zz_invSub_15 = invSboxRom_220;
      8'b11011101 : _zz_invSub_15 = invSboxRom_221;
      8'b11011110 : _zz_invSub_15 = invSboxRom_222;
      8'b11011111 : _zz_invSub_15 = invSboxRom_223;
      8'b11100000 : _zz_invSub_15 = invSboxRom_224;
      8'b11100001 : _zz_invSub_15 = invSboxRom_225;
      8'b11100010 : _zz_invSub_15 = invSboxRom_226;
      8'b11100011 : _zz_invSub_15 = invSboxRom_227;
      8'b11100100 : _zz_invSub_15 = invSboxRom_228;
      8'b11100101 : _zz_invSub_15 = invSboxRom_229;
      8'b11100110 : _zz_invSub_15 = invSboxRom_230;
      8'b11100111 : _zz_invSub_15 = invSboxRom_231;
      8'b11101000 : _zz_invSub_15 = invSboxRom_232;
      8'b11101001 : _zz_invSub_15 = invSboxRom_233;
      8'b11101010 : _zz_invSub_15 = invSboxRom_234;
      8'b11101011 : _zz_invSub_15 = invSboxRom_235;
      8'b11101100 : _zz_invSub_15 = invSboxRom_236;
      8'b11101101 : _zz_invSub_15 = invSboxRom_237;
      8'b11101110 : _zz_invSub_15 = invSboxRom_238;
      8'b11101111 : _zz_invSub_15 = invSboxRom_239;
      8'b11110000 : _zz_invSub_15 = invSboxRom_240;
      8'b11110001 : _zz_invSub_15 = invSboxRom_241;
      8'b11110010 : _zz_invSub_15 = invSboxRom_242;
      8'b11110011 : _zz_invSub_15 = invSboxRom_243;
      8'b11110100 : _zz_invSub_15 = invSboxRom_244;
      8'b11110101 : _zz_invSub_15 = invSboxRom_245;
      8'b11110110 : _zz_invSub_15 = invSboxRom_246;
      8'b11110111 : _zz_invSub_15 = invSboxRom_247;
      8'b11111000 : _zz_invSub_15 = invSboxRom_248;
      8'b11111001 : _zz_invSub_15 = invSboxRom_249;
      8'b11111010 : _zz_invSub_15 = invSboxRom_250;
      8'b11111011 : _zz_invSub_15 = invSboxRom_251;
      8'b11111100 : _zz_invSub_15 = invSboxRom_252;
      8'b11111101 : _zz_invSub_15 = invSboxRom_253;
      8'b11111110 : _zz_invSub_15 = invSboxRom_254;
      default : _zz_invSub_15 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_5_1)
      8'b00000000 : _zz__zz_roundKeyReg_0_5 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_5 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_5 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_5 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_5 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_5 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_5 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_5 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_5 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_5 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_5 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_5 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_5 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_5 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_5 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_5 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_5 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_5 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_5 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_5 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_5 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_5 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_5 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_5 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_5 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_5 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_5 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_5 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_5 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_5 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_5 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_5 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_5 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_5 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_5 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_5 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_5 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_5 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_5 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_5 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_5 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_5 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_5 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_5 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_5 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_5 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_5 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_5 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_5 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_5 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_5 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_5 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_5 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_5 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_5 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_5 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_5 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_5 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_5 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_5 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_5 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_5 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_5 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_5 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_5 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_5 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_5 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_5 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_5 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_5 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_5 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_5 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_5 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_5 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_5 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_5 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_5 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_5 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_5 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_5 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_5 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_5 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_5 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_5 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_5 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_5 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_5 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_5 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_5 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_5 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_5 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_5 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_5 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_5 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_5 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_5 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_5 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_5 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_5 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_5 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_5 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_5 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_5 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_5 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_5 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_5 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_5 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_5 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_5 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_5 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_5 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_5 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_5 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_5 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_5 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_5 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_5 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_5 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_5 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_5 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_5 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_5 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_5 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_5 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_5 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_5 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_5 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_5 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_5 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_5 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_5 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_5 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_5 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_5 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_5 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_5 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_5 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_5 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_5 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_5 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_5 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_5 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_5 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_5 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_5 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_5 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_5 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_5 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_5 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_5 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_5 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_5 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_5 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_5 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_5 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_5 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_5 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_5 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_5 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_5 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_5 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_5 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_5 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_5 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_5 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_5 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_5 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_5 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_5 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_5 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_5 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_5 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_5 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_5 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_5 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_5 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_5 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_5 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_5 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_5 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_5 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_5 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_5 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_5 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_5 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_5 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_5 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_5 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_5 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_5 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_5 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_5 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_5 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_5 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_5 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_5 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_5 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_5 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_5 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_5 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_5 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_5 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_5 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_5 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_5 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_5 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_5 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_5 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_5 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_5 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_5 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_5 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_5 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_5 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_5 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_5 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_5 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_5 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_5 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_5 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_5 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_5 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_5 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_5 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_5 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_5 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_5 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_5 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_5 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_5 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_5 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_5 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_5 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_5 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_5 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_5 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_5 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_5 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_5 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_5 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_5 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_5 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_5 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_5 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_5 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_5 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_5 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_5 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_5 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_5 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_5 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_5 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_5 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_5 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_5 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_5 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_5_3)
      8'b00000000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_5_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_5_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_5_5)
      8'b00000000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_5_4 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_5_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_5_7)
      8'b00000000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_5_6 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_5_6 = sboxRom_255;
    endcase
  end

  assign sboxRom_0 = 8'h63;
  assign sboxRom_1 = 8'h7c;
  assign sboxRom_2 = 8'h77;
  assign sboxRom_3 = 8'h7b;
  assign sboxRom_4 = 8'hf2;
  assign sboxRom_5 = 8'h6b;
  assign sboxRom_6 = 8'h6f;
  assign sboxRom_7 = 8'hc5;
  assign sboxRom_8 = 8'h30;
  assign sboxRom_9 = 8'h01;
  assign sboxRom_10 = 8'h67;
  assign sboxRom_11 = 8'h2b;
  assign sboxRom_12 = 8'hfe;
  assign sboxRom_13 = 8'hd7;
  assign sboxRom_14 = 8'hab;
  assign sboxRom_15 = 8'h76;
  assign sboxRom_16 = 8'hca;
  assign sboxRom_17 = 8'h82;
  assign sboxRom_18 = 8'hc9;
  assign sboxRom_19 = 8'h7d;
  assign sboxRom_20 = 8'hfa;
  assign sboxRom_21 = 8'h59;
  assign sboxRom_22 = 8'h47;
  assign sboxRom_23 = 8'hf0;
  assign sboxRom_24 = 8'had;
  assign sboxRom_25 = 8'hd4;
  assign sboxRom_26 = 8'ha2;
  assign sboxRom_27 = 8'haf;
  assign sboxRom_28 = 8'h9c;
  assign sboxRom_29 = 8'ha4;
  assign sboxRom_30 = 8'h72;
  assign sboxRom_31 = 8'hc0;
  assign sboxRom_32 = 8'hb7;
  assign sboxRom_33 = 8'hfd;
  assign sboxRom_34 = 8'h93;
  assign sboxRom_35 = 8'h26;
  assign sboxRom_36 = 8'h36;
  assign sboxRom_37 = 8'h3f;
  assign sboxRom_38 = 8'hf7;
  assign sboxRom_39 = 8'hcc;
  assign sboxRom_40 = 8'h34;
  assign sboxRom_41 = 8'ha5;
  assign sboxRom_42 = 8'he5;
  assign sboxRom_43 = 8'hf1;
  assign sboxRom_44 = 8'h71;
  assign sboxRom_45 = 8'hd8;
  assign sboxRom_46 = 8'h31;
  assign sboxRom_47 = 8'h15;
  assign sboxRom_48 = 8'h04;
  assign sboxRom_49 = 8'hc7;
  assign sboxRom_50 = 8'h23;
  assign sboxRom_51 = 8'hc3;
  assign sboxRom_52 = 8'h18;
  assign sboxRom_53 = 8'h96;
  assign sboxRom_54 = 8'h05;
  assign sboxRom_55 = 8'h9a;
  assign sboxRom_56 = 8'h07;
  assign sboxRom_57 = 8'h12;
  assign sboxRom_58 = 8'h80;
  assign sboxRom_59 = 8'he2;
  assign sboxRom_60 = 8'heb;
  assign sboxRom_61 = 8'h27;
  assign sboxRom_62 = 8'hb2;
  assign sboxRom_63 = 8'h75;
  assign sboxRom_64 = 8'h09;
  assign sboxRom_65 = 8'h83;
  assign sboxRom_66 = 8'h2c;
  assign sboxRom_67 = 8'h1a;
  assign sboxRom_68 = 8'h1b;
  assign sboxRom_69 = 8'h6e;
  assign sboxRom_70 = 8'h5a;
  assign sboxRom_71 = 8'ha0;
  assign sboxRom_72 = 8'h52;
  assign sboxRom_73 = 8'h3b;
  assign sboxRom_74 = 8'hd6;
  assign sboxRom_75 = 8'hb3;
  assign sboxRom_76 = 8'h29;
  assign sboxRom_77 = 8'he3;
  assign sboxRom_78 = 8'h2f;
  assign sboxRom_79 = 8'h84;
  assign sboxRom_80 = 8'h53;
  assign sboxRom_81 = 8'hd1;
  assign sboxRom_82 = 8'h0;
  assign sboxRom_83 = 8'hed;
  assign sboxRom_84 = 8'h20;
  assign sboxRom_85 = 8'hfc;
  assign sboxRom_86 = 8'hb1;
  assign sboxRom_87 = 8'h5b;
  assign sboxRom_88 = 8'h6a;
  assign sboxRom_89 = 8'hcb;
  assign sboxRom_90 = 8'hbe;
  assign sboxRom_91 = 8'h39;
  assign sboxRom_92 = 8'h4a;
  assign sboxRom_93 = 8'h4c;
  assign sboxRom_94 = 8'h58;
  assign sboxRom_95 = 8'hcf;
  assign sboxRom_96 = 8'hd0;
  assign sboxRom_97 = 8'hef;
  assign sboxRom_98 = 8'haa;
  assign sboxRom_99 = 8'hfb;
  assign sboxRom_100 = 8'h43;
  assign sboxRom_101 = 8'h4d;
  assign sboxRom_102 = 8'h33;
  assign sboxRom_103 = 8'h85;
  assign sboxRom_104 = 8'h45;
  assign sboxRom_105 = 8'hf9;
  assign sboxRom_106 = 8'h02;
  assign sboxRom_107 = 8'h7f;
  assign sboxRom_108 = 8'h50;
  assign sboxRom_109 = 8'h3c;
  assign sboxRom_110 = 8'h9f;
  assign sboxRom_111 = 8'ha8;
  assign sboxRom_112 = 8'h51;
  assign sboxRom_113 = 8'ha3;
  assign sboxRom_114 = 8'h40;
  assign sboxRom_115 = 8'h8f;
  assign sboxRom_116 = 8'h92;
  assign sboxRom_117 = 8'h9d;
  assign sboxRom_118 = 8'h38;
  assign sboxRom_119 = 8'hf5;
  assign sboxRom_120 = 8'hbc;
  assign sboxRom_121 = 8'hb6;
  assign sboxRom_122 = 8'hda;
  assign sboxRom_123 = 8'h21;
  assign sboxRom_124 = 8'h10;
  assign sboxRom_125 = 8'hff;
  assign sboxRom_126 = 8'hf3;
  assign sboxRom_127 = 8'hd2;
  assign sboxRom_128 = 8'hcd;
  assign sboxRom_129 = 8'h0c;
  assign sboxRom_130 = 8'h13;
  assign sboxRom_131 = 8'hec;
  assign sboxRom_132 = 8'h5f;
  assign sboxRom_133 = 8'h97;
  assign sboxRom_134 = 8'h44;
  assign sboxRom_135 = 8'h17;
  assign sboxRom_136 = 8'hc4;
  assign sboxRom_137 = 8'ha7;
  assign sboxRom_138 = 8'h7e;
  assign sboxRom_139 = 8'h3d;
  assign sboxRom_140 = 8'h64;
  assign sboxRom_141 = 8'h5d;
  assign sboxRom_142 = 8'h19;
  assign sboxRom_143 = 8'h73;
  assign sboxRom_144 = 8'h60;
  assign sboxRom_145 = 8'h81;
  assign sboxRom_146 = 8'h4f;
  assign sboxRom_147 = 8'hdc;
  assign sboxRom_148 = 8'h22;
  assign sboxRom_149 = 8'h2a;
  assign sboxRom_150 = 8'h90;
  assign sboxRom_151 = 8'h88;
  assign sboxRom_152 = 8'h46;
  assign sboxRom_153 = 8'hee;
  assign sboxRom_154 = 8'hb8;
  assign sboxRom_155 = 8'h14;
  assign sboxRom_156 = 8'hde;
  assign sboxRom_157 = 8'h5e;
  assign sboxRom_158 = 8'h0b;
  assign sboxRom_159 = 8'hdb;
  assign sboxRom_160 = 8'he0;
  assign sboxRom_161 = 8'h32;
  assign sboxRom_162 = 8'h3a;
  assign sboxRom_163 = 8'h0a;
  assign sboxRom_164 = 8'h49;
  assign sboxRom_165 = 8'h06;
  assign sboxRom_166 = 8'h24;
  assign sboxRom_167 = 8'h5c;
  assign sboxRom_168 = 8'hc2;
  assign sboxRom_169 = 8'hd3;
  assign sboxRom_170 = 8'hac;
  assign sboxRom_171 = 8'h62;
  assign sboxRom_172 = 8'h91;
  assign sboxRom_173 = 8'h95;
  assign sboxRom_174 = 8'he4;
  assign sboxRom_175 = 8'h79;
  assign sboxRom_176 = 8'he7;
  assign sboxRom_177 = 8'hc8;
  assign sboxRom_178 = 8'h37;
  assign sboxRom_179 = 8'h6d;
  assign sboxRom_180 = 8'h8d;
  assign sboxRom_181 = 8'hd5;
  assign sboxRom_182 = 8'h4e;
  assign sboxRom_183 = 8'ha9;
  assign sboxRom_184 = 8'h6c;
  assign sboxRom_185 = 8'h56;
  assign sboxRom_186 = 8'hf4;
  assign sboxRom_187 = 8'hea;
  assign sboxRom_188 = 8'h65;
  assign sboxRom_189 = 8'h7a;
  assign sboxRom_190 = 8'hae;
  assign sboxRom_191 = 8'h08;
  assign sboxRom_192 = 8'hba;
  assign sboxRom_193 = 8'h78;
  assign sboxRom_194 = 8'h25;
  assign sboxRom_195 = 8'h2e;
  assign sboxRom_196 = 8'h1c;
  assign sboxRom_197 = 8'ha6;
  assign sboxRom_198 = 8'hb4;
  assign sboxRom_199 = 8'hc6;
  assign sboxRom_200 = 8'he8;
  assign sboxRom_201 = 8'hdd;
  assign sboxRom_202 = 8'h74;
  assign sboxRom_203 = 8'h1f;
  assign sboxRom_204 = 8'h4b;
  assign sboxRom_205 = 8'hbd;
  assign sboxRom_206 = 8'h8b;
  assign sboxRom_207 = 8'h8a;
  assign sboxRom_208 = 8'h70;
  assign sboxRom_209 = 8'h3e;
  assign sboxRom_210 = 8'hb5;
  assign sboxRom_211 = 8'h66;
  assign sboxRom_212 = 8'h48;
  assign sboxRom_213 = 8'h03;
  assign sboxRom_214 = 8'hf6;
  assign sboxRom_215 = 8'h0e;
  assign sboxRom_216 = 8'h61;
  assign sboxRom_217 = 8'h35;
  assign sboxRom_218 = 8'h57;
  assign sboxRom_219 = 8'hb9;
  assign sboxRom_220 = 8'h86;
  assign sboxRom_221 = 8'hc1;
  assign sboxRom_222 = 8'h1d;
  assign sboxRom_223 = 8'h9e;
  assign sboxRom_224 = 8'he1;
  assign sboxRom_225 = 8'hf8;
  assign sboxRom_226 = 8'h98;
  assign sboxRom_227 = 8'h11;
  assign sboxRom_228 = 8'h69;
  assign sboxRom_229 = 8'hd9;
  assign sboxRom_230 = 8'h8e;
  assign sboxRom_231 = 8'h94;
  assign sboxRom_232 = 8'h9b;
  assign sboxRom_233 = 8'h1e;
  assign sboxRom_234 = 8'h87;
  assign sboxRom_235 = 8'he9;
  assign sboxRom_236 = 8'hce;
  assign sboxRom_237 = 8'h55;
  assign sboxRom_238 = 8'h28;
  assign sboxRom_239 = 8'hdf;
  assign sboxRom_240 = 8'h8c;
  assign sboxRom_241 = 8'ha1;
  assign sboxRom_242 = 8'h89;
  assign sboxRom_243 = 8'h0d;
  assign sboxRom_244 = 8'hbf;
  assign sboxRom_245 = 8'he6;
  assign sboxRom_246 = 8'h42;
  assign sboxRom_247 = 8'h68;
  assign sboxRom_248 = 8'h41;
  assign sboxRom_249 = 8'h99;
  assign sboxRom_250 = 8'h2d;
  assign sboxRom_251 = 8'h0f;
  assign sboxRom_252 = 8'hb0;
  assign sboxRom_253 = 8'h54;
  assign sboxRom_254 = 8'hbb;
  assign sboxRom_255 = 8'h16;
  assign rcon_0 = 8'h01;
  assign rcon_1 = 8'h02;
  assign rcon_2 = 8'h04;
  assign rcon_3 = 8'h08;
  assign rcon_4 = 8'h10;
  assign rcon_5 = 8'h20;
  assign rcon_6 = 8'h40;
  assign rcon_7 = 8'h80;
  assign rcon_8 = 8'h1b;
  assign rcon_9 = 8'h36;
  assign io_busy = running;
  always @(*) begin
    io_done = 1'b0;
    if(!when_AES128_l230) begin
      if(when_AES128_l244) begin
        if(when_AES128_l307) begin
          io_done = 1'b1;
        end
      end else begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              if(when_AES128_l397) begin
                io_done = 1'b1;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    io_dataOut = stateReg;
    if(!when_AES128_l230) begin
      if(when_AES128_l244) begin
        if(when_AES128_l307) begin
          io_dataOut = stateReg;
        end
      end else begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              if(when_AES128_l397) begin
                io_dataOut = stateReg;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    newStateComb = 128'h0;
    if(!when_AES128_l230) begin
      if(when_AES128_l244) begin
        newStateComb = _zz_stateReg_68;
      end
    end
  end

  always @(*) begin
    rkBitsUsedComb = 128'h0;
    if(!when_AES128_l230) begin
      if(when_AES128_l244) begin
        rkBitsUsedComb = _zz_stateReg_69;
      end
    end
  end

  assign invSboxRom_0 = 8'h52;
  assign invSboxRom_1 = 8'h09;
  assign invSboxRom_2 = 8'h6a;
  assign invSboxRom_3 = 8'hd5;
  assign invSboxRom_4 = 8'h30;
  assign invSboxRom_5 = 8'h36;
  assign invSboxRom_6 = 8'ha5;
  assign invSboxRom_7 = 8'h38;
  assign invSboxRom_8 = 8'hbf;
  assign invSboxRom_9 = 8'h40;
  assign invSboxRom_10 = 8'ha3;
  assign invSboxRom_11 = 8'h9e;
  assign invSboxRom_12 = 8'h81;
  assign invSboxRom_13 = 8'hf3;
  assign invSboxRom_14 = 8'hd7;
  assign invSboxRom_15 = 8'hfb;
  assign invSboxRom_16 = 8'h7c;
  assign invSboxRom_17 = 8'he3;
  assign invSboxRom_18 = 8'h39;
  assign invSboxRom_19 = 8'h82;
  assign invSboxRom_20 = 8'h9b;
  assign invSboxRom_21 = 8'h2f;
  assign invSboxRom_22 = 8'hff;
  assign invSboxRom_23 = 8'h87;
  assign invSboxRom_24 = 8'h34;
  assign invSboxRom_25 = 8'h8e;
  assign invSboxRom_26 = 8'h43;
  assign invSboxRom_27 = 8'h44;
  assign invSboxRom_28 = 8'hc4;
  assign invSboxRom_29 = 8'hde;
  assign invSboxRom_30 = 8'he9;
  assign invSboxRom_31 = 8'hcb;
  assign invSboxRom_32 = 8'h54;
  assign invSboxRom_33 = 8'h7b;
  assign invSboxRom_34 = 8'h94;
  assign invSboxRom_35 = 8'h32;
  assign invSboxRom_36 = 8'ha6;
  assign invSboxRom_37 = 8'hc2;
  assign invSboxRom_38 = 8'h23;
  assign invSboxRom_39 = 8'h3d;
  assign invSboxRom_40 = 8'hee;
  assign invSboxRom_41 = 8'h4c;
  assign invSboxRom_42 = 8'h95;
  assign invSboxRom_43 = 8'h0b;
  assign invSboxRom_44 = 8'h42;
  assign invSboxRom_45 = 8'hfa;
  assign invSboxRom_46 = 8'hc3;
  assign invSboxRom_47 = 8'h4e;
  assign invSboxRom_48 = 8'h08;
  assign invSboxRom_49 = 8'h2e;
  assign invSboxRom_50 = 8'ha1;
  assign invSboxRom_51 = 8'h66;
  assign invSboxRom_52 = 8'h28;
  assign invSboxRom_53 = 8'hd9;
  assign invSboxRom_54 = 8'h24;
  assign invSboxRom_55 = 8'hb2;
  assign invSboxRom_56 = 8'h76;
  assign invSboxRom_57 = 8'h5b;
  assign invSboxRom_58 = 8'ha2;
  assign invSboxRom_59 = 8'h49;
  assign invSboxRom_60 = 8'h6d;
  assign invSboxRom_61 = 8'h8b;
  assign invSboxRom_62 = 8'hd1;
  assign invSboxRom_63 = 8'h25;
  assign invSboxRom_64 = 8'h72;
  assign invSboxRom_65 = 8'hf8;
  assign invSboxRom_66 = 8'hf6;
  assign invSboxRom_67 = 8'h64;
  assign invSboxRom_68 = 8'h86;
  assign invSboxRom_69 = 8'h68;
  assign invSboxRom_70 = 8'h98;
  assign invSboxRom_71 = 8'h16;
  assign invSboxRom_72 = 8'hd4;
  assign invSboxRom_73 = 8'ha4;
  assign invSboxRom_74 = 8'h5c;
  assign invSboxRom_75 = 8'hcc;
  assign invSboxRom_76 = 8'h5d;
  assign invSboxRom_77 = 8'h65;
  assign invSboxRom_78 = 8'hb6;
  assign invSboxRom_79 = 8'h92;
  assign invSboxRom_80 = 8'h6c;
  assign invSboxRom_81 = 8'h70;
  assign invSboxRom_82 = 8'h48;
  assign invSboxRom_83 = 8'h50;
  assign invSboxRom_84 = 8'hfd;
  assign invSboxRom_85 = 8'hed;
  assign invSboxRom_86 = 8'hb9;
  assign invSboxRom_87 = 8'hda;
  assign invSboxRom_88 = 8'h5e;
  assign invSboxRom_89 = 8'h15;
  assign invSboxRom_90 = 8'h46;
  assign invSboxRom_91 = 8'h57;
  assign invSboxRom_92 = 8'ha7;
  assign invSboxRom_93 = 8'h8d;
  assign invSboxRom_94 = 8'h9d;
  assign invSboxRom_95 = 8'h84;
  assign invSboxRom_96 = 8'h90;
  assign invSboxRom_97 = 8'hd8;
  assign invSboxRom_98 = 8'hab;
  assign invSboxRom_99 = 8'h0;
  assign invSboxRom_100 = 8'h8c;
  assign invSboxRom_101 = 8'hbc;
  assign invSboxRom_102 = 8'hd3;
  assign invSboxRom_103 = 8'h0a;
  assign invSboxRom_104 = 8'hf7;
  assign invSboxRom_105 = 8'he4;
  assign invSboxRom_106 = 8'h58;
  assign invSboxRom_107 = 8'h05;
  assign invSboxRom_108 = 8'hb8;
  assign invSboxRom_109 = 8'hb3;
  assign invSboxRom_110 = 8'h45;
  assign invSboxRom_111 = 8'h06;
  assign invSboxRom_112 = 8'hd0;
  assign invSboxRom_113 = 8'h2c;
  assign invSboxRom_114 = 8'h1e;
  assign invSboxRom_115 = 8'h8f;
  assign invSboxRom_116 = 8'hca;
  assign invSboxRom_117 = 8'h3f;
  assign invSboxRom_118 = 8'h0f;
  assign invSboxRom_119 = 8'h02;
  assign invSboxRom_120 = 8'hc1;
  assign invSboxRom_121 = 8'haf;
  assign invSboxRom_122 = 8'hbd;
  assign invSboxRom_123 = 8'h03;
  assign invSboxRom_124 = 8'h01;
  assign invSboxRom_125 = 8'h13;
  assign invSboxRom_126 = 8'h8a;
  assign invSboxRom_127 = 8'h6b;
  assign invSboxRom_128 = 8'h3a;
  assign invSboxRom_129 = 8'h91;
  assign invSboxRom_130 = 8'h11;
  assign invSboxRom_131 = 8'h41;
  assign invSboxRom_132 = 8'h4f;
  assign invSboxRom_133 = 8'h67;
  assign invSboxRom_134 = 8'hdc;
  assign invSboxRom_135 = 8'hea;
  assign invSboxRom_136 = 8'h97;
  assign invSboxRom_137 = 8'hf2;
  assign invSboxRom_138 = 8'hcf;
  assign invSboxRom_139 = 8'hce;
  assign invSboxRom_140 = 8'hf0;
  assign invSboxRom_141 = 8'hb4;
  assign invSboxRom_142 = 8'he6;
  assign invSboxRom_143 = 8'h73;
  assign invSboxRom_144 = 8'h96;
  assign invSboxRom_145 = 8'hac;
  assign invSboxRom_146 = 8'h74;
  assign invSboxRom_147 = 8'h22;
  assign invSboxRom_148 = 8'he7;
  assign invSboxRom_149 = 8'had;
  assign invSboxRom_150 = 8'h35;
  assign invSboxRom_151 = 8'h85;
  assign invSboxRom_152 = 8'he2;
  assign invSboxRom_153 = 8'hf9;
  assign invSboxRom_154 = 8'h37;
  assign invSboxRom_155 = 8'he8;
  assign invSboxRom_156 = 8'h1c;
  assign invSboxRom_157 = 8'h75;
  assign invSboxRom_158 = 8'hdf;
  assign invSboxRom_159 = 8'h6e;
  assign invSboxRom_160 = 8'h47;
  assign invSboxRom_161 = 8'hf1;
  assign invSboxRom_162 = 8'h1a;
  assign invSboxRom_163 = 8'h71;
  assign invSboxRom_164 = 8'h1d;
  assign invSboxRom_165 = 8'h29;
  assign invSboxRom_166 = 8'hc5;
  assign invSboxRom_167 = 8'h89;
  assign invSboxRom_168 = 8'h6f;
  assign invSboxRom_169 = 8'hb7;
  assign invSboxRom_170 = 8'h62;
  assign invSboxRom_171 = 8'h0e;
  assign invSboxRom_172 = 8'haa;
  assign invSboxRom_173 = 8'h18;
  assign invSboxRom_174 = 8'hbe;
  assign invSboxRom_175 = 8'h1b;
  assign invSboxRom_176 = 8'hfc;
  assign invSboxRom_177 = 8'h56;
  assign invSboxRom_178 = 8'h3e;
  assign invSboxRom_179 = 8'h4b;
  assign invSboxRom_180 = 8'hc6;
  assign invSboxRom_181 = 8'hd2;
  assign invSboxRom_182 = 8'h79;
  assign invSboxRom_183 = 8'h20;
  assign invSboxRom_184 = 8'h9a;
  assign invSboxRom_185 = 8'hdb;
  assign invSboxRom_186 = 8'hc0;
  assign invSboxRom_187 = 8'hfe;
  assign invSboxRom_188 = 8'h78;
  assign invSboxRom_189 = 8'hcd;
  assign invSboxRom_190 = 8'h5a;
  assign invSboxRom_191 = 8'hf4;
  assign invSboxRom_192 = 8'h1f;
  assign invSboxRom_193 = 8'hdd;
  assign invSboxRom_194 = 8'ha8;
  assign invSboxRom_195 = 8'h33;
  assign invSboxRom_196 = 8'h88;
  assign invSboxRom_197 = 8'h07;
  assign invSboxRom_198 = 8'hc7;
  assign invSboxRom_199 = 8'h31;
  assign invSboxRom_200 = 8'hb1;
  assign invSboxRom_201 = 8'h12;
  assign invSboxRom_202 = 8'h10;
  assign invSboxRom_203 = 8'h59;
  assign invSboxRom_204 = 8'h27;
  assign invSboxRom_205 = 8'h80;
  assign invSboxRom_206 = 8'hec;
  assign invSboxRom_207 = 8'h5f;
  assign invSboxRom_208 = 8'h60;
  assign invSboxRom_209 = 8'h51;
  assign invSboxRom_210 = 8'h7f;
  assign invSboxRom_211 = 8'ha9;
  assign invSboxRom_212 = 8'h19;
  assign invSboxRom_213 = 8'hb5;
  assign invSboxRom_214 = 8'h4a;
  assign invSboxRom_215 = 8'h0d;
  assign invSboxRom_216 = 8'h2d;
  assign invSboxRom_217 = 8'he5;
  assign invSboxRom_218 = 8'h7a;
  assign invSboxRom_219 = 8'h9f;
  assign invSboxRom_220 = 8'h93;
  assign invSboxRom_221 = 8'hc9;
  assign invSboxRom_222 = 8'h9c;
  assign invSboxRom_223 = 8'hef;
  assign invSboxRom_224 = 8'ha0;
  assign invSboxRom_225 = 8'he0;
  assign invSboxRom_226 = 8'h3b;
  assign invSboxRom_227 = 8'h4d;
  assign invSboxRom_228 = 8'hae;
  assign invSboxRom_229 = 8'h2a;
  assign invSboxRom_230 = 8'hf5;
  assign invSboxRom_231 = 8'hb0;
  assign invSboxRom_232 = 8'hc8;
  assign invSboxRom_233 = 8'heb;
  assign invSboxRom_234 = 8'hbb;
  assign invSboxRom_235 = 8'h3c;
  assign invSboxRom_236 = 8'h83;
  assign invSboxRom_237 = 8'h53;
  assign invSboxRom_238 = 8'h99;
  assign invSboxRom_239 = 8'h61;
  assign invSboxRom_240 = 8'h17;
  assign invSboxRom_241 = 8'h2b;
  assign invSboxRom_242 = 8'h04;
  assign invSboxRom_243 = 8'h7e;
  assign invSboxRom_244 = 8'hba;
  assign invSboxRom_245 = 8'h77;
  assign invSboxRom_246 = 8'hd6;
  assign invSboxRom_247 = 8'h26;
  assign invSboxRom_248 = 8'he1;
  assign invSboxRom_249 = 8'h69;
  assign invSboxRom_250 = 8'h14;
  assign invSboxRom_251 = 8'h63;
  assign invSboxRom_252 = 8'h55;
  assign invSboxRom_253 = 8'h21;
  assign invSboxRom_254 = 8'h0c;
  assign invSboxRom_255 = 8'h7d;
  always @(*) begin
    initKeyWords_0 = 32'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(when_AES128_l315) begin
          initKeyWords_0 = _zz_roundKeyReg_0_3;
        end
      end
    end
  end

  always @(*) begin
    initKeyWords_1 = 32'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(when_AES128_l315) begin
          initKeyWords_1 = _zz_roundKeyReg_1_1;
        end
      end
    end
  end

  always @(*) begin
    initKeyWords_2 = 32'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(when_AES128_l315) begin
          initKeyWords_2 = _zz_roundKeyReg_2_1;
        end
      end
    end
  end

  always @(*) begin
    initKeyWords_3 = 32'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(when_AES128_l315) begin
          initKeyWords_3 = _zz_roundKeyReg_3_1;
        end
      end
    end
  end

  always @(*) begin
    invShifted_0 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_0 = stateReg[127 : 120];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_0 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_0 = _zz_invSub_0;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_0 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_0 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_0 = _zz_invMixed_0_1;
              end else begin
                invMixed_0 = (((((_zz_invMixed_0_33 ^ _zz_invMixed_0_34) ^ (_zz_invMixed_0_35 ? _zz_invMixed_0_36 : _zz_invMixed_0_13)) ^ ((_zz_invMixed_0_37 ^ _zz_invMixed_0_38) ^ _zz_invMixed_0_2)) ^ (((_zz_invMixed_0_39 ? _zz_invMixed_0_40 : _zz_invMixed_0_24) ^ (_zz_invMixed_0_41 ? _zz_invMixed_0_42 : _zz_invMixed_0_27)) ^ _zz_invMixed_0_3)) ^ ((_zz_invMixed_0_31[7] ? (_zz_invMixed_0_32 ^ 8'h1b) : _zz_invMixed_0_32) ^ _zz_invMixed_0_4));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_1 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_1 = stateReg[23 : 16];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_1 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_1 = _zz_invSub_1;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_1 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_1 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_1 = _zz_invMixed_0_2;
              end else begin
                invMixed_1 = (((((_zz_invMixed_1_28 ? _zz_invMixed_1_29 : _zz_invMixed_1_4) ^ _zz_invMixed_0_1) ^ ((_zz_invMixed_1_30 ^ _zz_invMixed_1_31) ^ (_zz_invMixed_1_32 ? _zz_invMixed_1_33 : _zz_invMixed_1_13))) ^ (((_zz_invMixed_1_34 ? _zz_invMixed_1_35 : _zz_invMixed_1_18) ^ (_zz_invMixed_1_36 ? _zz_invMixed_1_37 : _zz_invMixed_1_19)) ^ _zz_invMixed_0_3)) ^ (((_zz_invMixed_1_23[7] ? (_zz_invMixed_1_24 ^ _zz_invMixed_1_38) : _zz_invMixed_1_24) ^ (_zz_invMixed_1_26[7] ? (_zz_invMixed_1_27 ^ _zz_invMixed_1_39) : _zz_invMixed_1_27)) ^ _zz_invMixed_0_4));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_2 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_2 = stateReg[47 : 40];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_2 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_2 = _zz_invSub_2;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_2 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_2 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_2 = _zz_invMixed_0_3;
              end else begin
                invMixed_2 = (((((_zz_invMixed_2_28 ^ _zz_invMixed_2_29) ^ _zz_invMixed_0_1) ^ ((_zz_invMixed_2_30 ? _zz_invMixed_2_31 : _zz_invMixed_2_12) ^ _zz_invMixed_0_2)) ^ (((_zz_invMixed_2_32 ? _zz_invMixed_2_33 : _zz_invMixed_2_17) ^ (_zz_invMixed_2_34 ? _zz_invMixed_2_35 : _zz_invMixed_2_20)) ^ (_zz_invMixed_0_3[7] ? (_zz_invMixed_2_21 ^ _zz_invMixed_2_36) : _zz_invMixed_2_21))) ^ (((_zz_invMixed_2_25[7] ? (_zz_invMixed_2_26 ^ _zz_invMixed_2_37) : _zz_invMixed_2_26) ^ (_zz_invMixed_0_4[7] ? (_zz_invMixed_2_27 ^ _zz_invMixed_2_38) : _zz_invMixed_2_27)) ^ _zz_invMixed_0_4));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_3 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_3 = stateReg[71 : 64];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_3 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_3 = _zz_invSub_3;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_3 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_3 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_3 = _zz_invMixed_0_4;
              end else begin
                invMixed_3 = (((((_zz_invMixed_3_28 ^ _zz_invMixed_3_29) ^ _zz_invMixed_0_1) ^ ((_zz_invMixed_3_30 ^ _zz_invMixed_3_31) ^ _zz_invMixed_0_2)) ^ ((_zz_invMixed_3_17[7] ? (_zz_invMixed_3_18 ^ _zz_invMixed_3_32) : _zz_invMixed_3_18) ^ _zz_invMixed_0_3)) ^ (((_zz_invMixed_3_22[7] ? (_zz_invMixed_3_23 ^ _zz_invMixed_3_33) : _zz_invMixed_3_23) ^ (_zz_invMixed_3_25[7] ? (_zz_invMixed_3_26 ^ _zz_invMixed_3_34) : _zz_invMixed_3_26)) ^ (_zz_invMixed_0_4[7] ? (_zz_invMixed_3_27 ^ 8'h1b) : _zz_invMixed_3_27)));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_4 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_4 = stateReg[95 : 88];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_4 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_4 = _zz_invSub_4;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_4 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_4 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_4 = _zz_invMixed_4;
              end else begin
                invMixed_4 = (((((_zz_invMixed_4_32 ^ _zz_invMixed_4_33) ^ (_zz_invMixed_4_34 ? _zz_invMixed_4_35 : _zz_invMixed_4_12)) ^ ((_zz_invMixed_4_36 ^ _zz_invMixed_4_37) ^ _zz_invMixed_4_1)) ^ (((_zz_invMixed_4_38 ? _zz_invMixed_4_39 : _zz_invMixed_4_23) ^ (_zz_invMixed_4_40 ? _zz_invMixed_4_41 : _zz_invMixed_4_26)) ^ _zz_invMixed_4_2)) ^ ((_zz_invMixed_4_30[7] ? (_zz_invMixed_4_31 ^ 8'h1b) : _zz_invMixed_4_31) ^ _zz_invMixed_4_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_5 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_5 = stateReg[119 : 112];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_5 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_5 = _zz_invSub_5;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_5 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_5 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_5 = _zz_invMixed_4_1;
              end else begin
                invMixed_5 = (((((_zz_invMixed_5_28 ? _zz_invMixed_5_29 : _zz_invMixed_5_4) ^ _zz_invMixed_4) ^ ((_zz_invMixed_5_30 ^ _zz_invMixed_5_31) ^ (_zz_invMixed_5_32 ? _zz_invMixed_5_33 : _zz_invMixed_5_13))) ^ (((_zz_invMixed_5_34 ? _zz_invMixed_5_35 : _zz_invMixed_5_18) ^ (_zz_invMixed_5_36 ? _zz_invMixed_5_37 : _zz_invMixed_5_19)) ^ _zz_invMixed_4_2)) ^ (((_zz_invMixed_5_23[7] ? (_zz_invMixed_5_24 ^ _zz_invMixed_5_38) : _zz_invMixed_5_24) ^ (_zz_invMixed_5_26[7] ? (_zz_invMixed_5_27 ^ _zz_invMixed_5_39) : _zz_invMixed_5_27)) ^ _zz_invMixed_4_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_6 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_6 = stateReg[15 : 8];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_6 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_6 = _zz_invSub_6;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_6 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_6 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_6 = _zz_invMixed_4_2;
              end else begin
                invMixed_6 = (((((_zz_invMixed_6_28 ^ _zz_invMixed_6_29) ^ _zz_invMixed_4) ^ ((_zz_invMixed_6_30 ? _zz_invMixed_6_31 : _zz_invMixed_6_12) ^ _zz_invMixed_4_1)) ^ (((_zz_invMixed_6_32 ? _zz_invMixed_6_33 : _zz_invMixed_6_17) ^ (_zz_invMixed_6_34 ? _zz_invMixed_6_35 : _zz_invMixed_6_20)) ^ (_zz_invMixed_4_2[7] ? (_zz_invMixed_6_21 ^ _zz_invMixed_6_36) : _zz_invMixed_6_21))) ^ (((_zz_invMixed_6_25[7] ? (_zz_invMixed_6_26 ^ _zz_invMixed_6_37) : _zz_invMixed_6_26) ^ (_zz_invMixed_4_3[7] ? (_zz_invMixed_6_27 ^ _zz_invMixed_6_38) : _zz_invMixed_6_27)) ^ _zz_invMixed_4_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_7 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_7 = stateReg[39 : 32];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_7 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_7 = _zz_invSub_7;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_7 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_7 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_7 = _zz_invMixed_4_3;
              end else begin
                invMixed_7 = (((((_zz_invMixed_7_28 ^ _zz_invMixed_7_29) ^ _zz_invMixed_4) ^ ((_zz_invMixed_7_30 ^ _zz_invMixed_7_31) ^ _zz_invMixed_4_1)) ^ ((_zz_invMixed_7_17[7] ? (_zz_invMixed_7_18 ^ _zz_invMixed_7_32) : _zz_invMixed_7_18) ^ _zz_invMixed_4_2)) ^ (((_zz_invMixed_7_22[7] ? (_zz_invMixed_7_23 ^ _zz_invMixed_7_33) : _zz_invMixed_7_23) ^ (_zz_invMixed_7_25[7] ? (_zz_invMixed_7_26 ^ _zz_invMixed_7_34) : _zz_invMixed_7_26)) ^ (_zz_invMixed_4_3[7] ? (_zz_invMixed_7_27 ^ 8'h1b) : _zz_invMixed_7_27)));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_8 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_8 = stateReg[63 : 56];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_8 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_8 = _zz_invSub_8;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_8 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_8 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_8 = _zz_invMixed_8;
              end else begin
                invMixed_8 = (((((_zz_invMixed_8_32 ^ _zz_invMixed_8_33) ^ (_zz_invMixed_8_34 ? _zz_invMixed_8_35 : _zz_invMixed_8_12)) ^ ((_zz_invMixed_8_36 ^ _zz_invMixed_8_37) ^ _zz_invMixed_8_1)) ^ (((_zz_invMixed_8_38 ? _zz_invMixed_8_39 : _zz_invMixed_8_23) ^ (_zz_invMixed_8_40 ? _zz_invMixed_8_41 : _zz_invMixed_8_26)) ^ _zz_invMixed_8_2)) ^ ((_zz_invMixed_8_30[7] ? (_zz_invMixed_8_31 ^ 8'h1b) : _zz_invMixed_8_31) ^ _zz_invMixed_8_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_9 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_9 = stateReg[87 : 80];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_9 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_9 = _zz_invSub_9;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_9 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_9 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_9 = _zz_invMixed_8_1;
              end else begin
                invMixed_9 = (((((_zz_invMixed_9_28 ? _zz_invMixed_9_29 : _zz_invMixed_9_4) ^ _zz_invMixed_8) ^ ((_zz_invMixed_9_30 ^ _zz_invMixed_9_31) ^ (_zz_invMixed_9_32 ? _zz_invMixed_9_33 : _zz_invMixed_9_13))) ^ (((_zz_invMixed_9_34 ? _zz_invMixed_9_35 : _zz_invMixed_9_18) ^ (_zz_invMixed_9_36 ? _zz_invMixed_9_37 : _zz_invMixed_9_19)) ^ _zz_invMixed_8_2)) ^ (((_zz_invMixed_9_23[7] ? (_zz_invMixed_9_24 ^ _zz_invMixed_9_38) : _zz_invMixed_9_24) ^ (_zz_invMixed_9_26[7] ? (_zz_invMixed_9_27 ^ _zz_invMixed_9_39) : _zz_invMixed_9_27)) ^ _zz_invMixed_8_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_10 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_10 = stateReg[111 : 104];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_10 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_10 = _zz_invSub_10;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_10 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_10 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_10 = _zz_invMixed_8_2;
              end else begin
                invMixed_10 = (((((_zz_invMixed_10_28 ^ _zz_invMixed_10_29) ^ _zz_invMixed_8) ^ ((_zz_invMixed_10_30 ? _zz_invMixed_10_31 : _zz_invMixed_10_12) ^ _zz_invMixed_8_1)) ^ (((_zz_invMixed_10_32 ? _zz_invMixed_10_33 : _zz_invMixed_10_17) ^ (_zz_invMixed_10_34 ? _zz_invMixed_10_35 : _zz_invMixed_10_20)) ^ (_zz_invMixed_8_2[7] ? (_zz_invMixed_10_21 ^ _zz_invMixed_10_36) : _zz_invMixed_10_21))) ^ (((_zz_invMixed_10_25[7] ? (_zz_invMixed_10_26 ^ _zz_invMixed_10_37) : _zz_invMixed_10_26) ^ (_zz_invMixed_8_3[7] ? (_zz_invMixed_10_27 ^ _zz_invMixed_10_38) : _zz_invMixed_10_27)) ^ _zz_invMixed_8_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_11 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_11 = stateReg[7 : 0];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_11 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_11 = _zz_invSub_11;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_11 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_11 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_11 = _zz_invMixed_8_3;
              end else begin
                invMixed_11 = (((((_zz_invMixed_11_28 ^ _zz_invMixed_11_29) ^ _zz_invMixed_8) ^ ((_zz_invMixed_11_30 ^ _zz_invMixed_11_31) ^ _zz_invMixed_8_1)) ^ ((_zz_invMixed_11_17[7] ? (_zz_invMixed_11_18 ^ _zz_invMixed_11_32) : _zz_invMixed_11_18) ^ _zz_invMixed_8_2)) ^ (((_zz_invMixed_11_22[7] ? (_zz_invMixed_11_23 ^ _zz_invMixed_11_33) : _zz_invMixed_11_23) ^ (_zz_invMixed_11_25[7] ? (_zz_invMixed_11_26 ^ _zz_invMixed_11_34) : _zz_invMixed_11_26)) ^ (_zz_invMixed_8_3[7] ? (_zz_invMixed_11_27 ^ 8'h1b) : _zz_invMixed_11_27)));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_12 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_12 = stateReg[31 : 24];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_12 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_12 = _zz_invSub_12;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_12 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_12 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_12 = _zz_invMixed_12;
              end else begin
                invMixed_12 = (((((_zz_invMixed_12_32 ^ _zz_invMixed_12_33) ^ (_zz_invMixed_12_34 ? _zz_invMixed_12_35 : _zz_invMixed_12_12)) ^ ((_zz_invMixed_12_36 ^ _zz_invMixed_12_37) ^ _zz_invMixed_12_1)) ^ (((_zz_invMixed_12_38 ? _zz_invMixed_12_39 : _zz_invMixed_12_23) ^ (_zz_invMixed_12_40 ? _zz_invMixed_12_41 : _zz_invMixed_12_26)) ^ _zz_invMixed_12_2)) ^ ((_zz_invMixed_12_30[7] ? (_zz_invMixed_12_31 ^ 8'h1b) : _zz_invMixed_12_31) ^ _zz_invMixed_12_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_13 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_13 = stateReg[55 : 48];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_13 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_13 = _zz_invSub_13;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_13 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_13 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_13 = _zz_invMixed_12_1;
              end else begin
                invMixed_13 = (((((_zz_invMixed_13_28 ? _zz_invMixed_13_29 : _zz_invMixed_13_4) ^ _zz_invMixed_12) ^ ((_zz_invMixed_13_30 ^ _zz_invMixed_13_31) ^ (_zz_invMixed_13_32 ? _zz_invMixed_13_33 : _zz_invMixed_13_13))) ^ (((_zz_invMixed_13_34 ? _zz_invMixed_13_35 : _zz_invMixed_13_18) ^ (_zz_invMixed_13_36 ? _zz_invMixed_13_37 : _zz_invMixed_13_19)) ^ _zz_invMixed_12_2)) ^ (((_zz_invMixed_13_23[7] ? (_zz_invMixed_13_24 ^ _zz_invMixed_13_38) : _zz_invMixed_13_24) ^ (_zz_invMixed_13_26[7] ? (_zz_invMixed_13_27 ^ _zz_invMixed_13_39) : _zz_invMixed_13_27)) ^ _zz_invMixed_12_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_14 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_14 = stateReg[79 : 72];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_14 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_14 = _zz_invSub_14;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_14 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_14 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_14 = _zz_invMixed_12_2;
              end else begin
                invMixed_14 = (((((_zz_invMixed_14_28 ^ _zz_invMixed_14_29) ^ _zz_invMixed_12) ^ ((_zz_invMixed_14_30 ? _zz_invMixed_14_31 : _zz_invMixed_14_12) ^ _zz_invMixed_12_1)) ^ (((_zz_invMixed_14_32 ? _zz_invMixed_14_33 : _zz_invMixed_14_17) ^ (_zz_invMixed_14_34 ? _zz_invMixed_14_35 : _zz_invMixed_14_20)) ^ (_zz_invMixed_12_2[7] ? (_zz_invMixed_14_21 ^ _zz_invMixed_14_36) : _zz_invMixed_14_21))) ^ (((_zz_invMixed_14_25[7] ? (_zz_invMixed_14_26 ^ _zz_invMixed_14_37) : _zz_invMixed_14_26) ^ (_zz_invMixed_12_3[7] ? (_zz_invMixed_14_27 ^ _zz_invMixed_14_38) : _zz_invMixed_14_27)) ^ _zz_invMixed_12_3));
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invShifted_15 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invShifted_15 = stateReg[103 : 96];
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invSub_15 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invSub_15 = _zz_invSub_15;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    invMixed_15 = 8'h0;
    if(!when_AES128_l230) begin
      if(!when_AES128_l244) begin
        if(!when_AES128_l315) begin
          if(!precomputeRunning) begin
            if(when_AES128_l339) begin
              invMixed_15 = 8'h0;
              if(when_AES128_l370) begin
                invMixed_15 = _zz_invMixed_12_3;
              end else begin
                invMixed_15 = (((((_zz_invMixed_15_28 ^ _zz_invMixed_15_29) ^ _zz_invMixed_12) ^ ((_zz_invMixed_15_30 ^ _zz_invMixed_15_31) ^ _zz_invMixed_12_1)) ^ ((_zz_invMixed_15_17[7] ? (_zz_invMixed_15_18 ^ _zz_invMixed_15_32) : _zz_invMixed_15_18) ^ _zz_invMixed_12_2)) ^ (((_zz_invMixed_15_22[7] ? (_zz_invMixed_15_23 ^ _zz_invMixed_15_33) : _zz_invMixed_15_23) ^ (_zz_invMixed_15_25[7] ? (_zz_invMixed_15_26 ^ _zz_invMixed_15_34) : _zz_invMixed_15_26)) ^ (_zz_invMixed_12_3[7] ? (_zz_invMixed_15_27 ^ 8'h1b) : _zz_invMixed_15_27)));
              end
            end
          end
        end
      end
    end
  end

  assign when_AES128_l230 = ((io_start && (! running)) && (! io_decrypt));
  assign _zz_stateReg = io_key[127 : 96];
  assign _zz_stateReg_1 = io_key[95 : 64];
  assign _zz_stateReg_2 = io_key[63 : 32];
  assign _zz_stateReg_3 = io_key[31 : 0];
  assign _zz_stateReg_4 = _zz__zz_stateReg_4;
  assign _zz_stateReg_8 = _zz__zz_stateReg_8;
  assign _zz_stateReg_12 = _zz__zz_stateReg_12;
  assign _zz_stateReg_16 = _zz__zz_stateReg_16;
  assign _zz_stateReg_5 = _zz__zz_stateReg_5;
  assign _zz_stateReg_9 = _zz__zz_stateReg_9;
  assign _zz_stateReg_13 = _zz__zz_stateReg_13;
  assign _zz_stateReg_17 = _zz__zz_stateReg_17;
  assign _zz_stateReg_6 = _zz__zz_stateReg_6;
  assign _zz_stateReg_10 = _zz__zz_stateReg_10;
  assign _zz_stateReg_14 = _zz__zz_stateReg_14;
  assign _zz_stateReg_18 = _zz__zz_stateReg_18;
  assign _zz_stateReg_7 = _zz__zz_stateReg_7;
  assign _zz_stateReg_11 = _zz__zz_stateReg_11;
  assign _zz_stateReg_15 = _zz__zz_stateReg_15;
  assign _zz_stateReg_19 = _zz__zz_stateReg_19;
  assign when_AES128_l272 = (roundCount == 4'b1001);
  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_20 = _zz_stateReg_4;
    end else begin
      _zz_stateReg_20 = ((((_zz_stateReg_4[7] ? (_zz_stateReg_36 ^ 8'h1b) : _zz_stateReg_36) ^ ((_zz_stateReg_5[7] ? (_zz_stateReg_37 ^ 8'h1b) : _zz_stateReg_37) ^ _zz_stateReg_5)) ^ _zz_stateReg_6) ^ _zz_stateReg_7);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_21 = _zz_stateReg_5;
    end else begin
      _zz_stateReg_21 = (((_zz_stateReg_4 ^ (_zz_stateReg_5[7] ? (_zz_stateReg_38 ^ 8'h1b) : _zz_stateReg_38)) ^ ((_zz_stateReg_6[7] ? (_zz_stateReg_39 ^ 8'h1b) : _zz_stateReg_39) ^ _zz_stateReg_6)) ^ _zz_stateReg_7);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_22 = _zz_stateReg_6;
    end else begin
      _zz_stateReg_22 = (((_zz_stateReg_4 ^ _zz_stateReg_5) ^ (_zz_stateReg_6[7] ? (_zz_stateReg_40 ^ 8'h1b) : _zz_stateReg_40)) ^ ((_zz_stateReg_7[7] ? (_zz_stateReg_41 ^ 8'h1b) : _zz_stateReg_41) ^ _zz_stateReg_7));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_23 = _zz_stateReg_7;
    end else begin
      _zz_stateReg_23 = (((((_zz_stateReg_4[7] ? (_zz_stateReg_42 ^ 8'h1b) : _zz_stateReg_42) ^ _zz_stateReg_4) ^ _zz_stateReg_5) ^ _zz_stateReg_6) ^ (_zz_stateReg_7[7] ? (_zz_stateReg_43 ^ 8'h1b) : _zz_stateReg_43));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_24 = _zz_stateReg_8;
    end else begin
      _zz_stateReg_24 = ((((_zz_stateReg_8[7] ? (_zz_stateReg_44 ^ 8'h1b) : _zz_stateReg_44) ^ ((_zz_stateReg_9[7] ? (_zz_stateReg_45 ^ 8'h1b) : _zz_stateReg_45) ^ _zz_stateReg_9)) ^ _zz_stateReg_10) ^ _zz_stateReg_11);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_25 = _zz_stateReg_9;
    end else begin
      _zz_stateReg_25 = (((_zz_stateReg_8 ^ (_zz_stateReg_9[7] ? (_zz_stateReg_46 ^ 8'h1b) : _zz_stateReg_46)) ^ ((_zz_stateReg_10[7] ? (_zz_stateReg_47 ^ 8'h1b) : _zz_stateReg_47) ^ _zz_stateReg_10)) ^ _zz_stateReg_11);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_26 = _zz_stateReg_10;
    end else begin
      _zz_stateReg_26 = (((_zz_stateReg_8 ^ _zz_stateReg_9) ^ (_zz_stateReg_10[7] ? (_zz_stateReg_48 ^ 8'h1b) : _zz_stateReg_48)) ^ ((_zz_stateReg_11[7] ? (_zz_stateReg_49 ^ 8'h1b) : _zz_stateReg_49) ^ _zz_stateReg_11));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_27 = _zz_stateReg_11;
    end else begin
      _zz_stateReg_27 = (((((_zz_stateReg_8[7] ? (_zz_stateReg_50 ^ 8'h1b) : _zz_stateReg_50) ^ _zz_stateReg_8) ^ _zz_stateReg_9) ^ _zz_stateReg_10) ^ (_zz_stateReg_11[7] ? (_zz_stateReg_51 ^ 8'h1b) : _zz_stateReg_51));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_28 = _zz_stateReg_12;
    end else begin
      _zz_stateReg_28 = ((((_zz_stateReg_12[7] ? (_zz_stateReg_52 ^ 8'h1b) : _zz_stateReg_52) ^ ((_zz_stateReg_13[7] ? (_zz_stateReg_53 ^ 8'h1b) : _zz_stateReg_53) ^ _zz_stateReg_13)) ^ _zz_stateReg_14) ^ _zz_stateReg_15);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_29 = _zz_stateReg_13;
    end else begin
      _zz_stateReg_29 = (((_zz_stateReg_12 ^ (_zz_stateReg_13[7] ? (_zz_stateReg_54 ^ 8'h1b) : _zz_stateReg_54)) ^ ((_zz_stateReg_14[7] ? (_zz_stateReg_55 ^ 8'h1b) : _zz_stateReg_55) ^ _zz_stateReg_14)) ^ _zz_stateReg_15);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_30 = _zz_stateReg_14;
    end else begin
      _zz_stateReg_30 = (((_zz_stateReg_12 ^ _zz_stateReg_13) ^ (_zz_stateReg_14[7] ? (_zz_stateReg_56 ^ 8'h1b) : _zz_stateReg_56)) ^ ((_zz_stateReg_15[7] ? (_zz_stateReg_57 ^ 8'h1b) : _zz_stateReg_57) ^ _zz_stateReg_15));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_31 = _zz_stateReg_15;
    end else begin
      _zz_stateReg_31 = (((((_zz_stateReg_12[7] ? (_zz_stateReg_58 ^ 8'h1b) : _zz_stateReg_58) ^ _zz_stateReg_12) ^ _zz_stateReg_13) ^ _zz_stateReg_14) ^ (_zz_stateReg_15[7] ? (_zz_stateReg_59 ^ 8'h1b) : _zz_stateReg_59));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_32 = _zz_stateReg_16;
    end else begin
      _zz_stateReg_32 = ((((_zz_stateReg_16[7] ? (_zz_stateReg_60 ^ 8'h1b) : _zz_stateReg_60) ^ ((_zz_stateReg_17[7] ? (_zz_stateReg_61 ^ 8'h1b) : _zz_stateReg_61) ^ _zz_stateReg_17)) ^ _zz_stateReg_18) ^ _zz_stateReg_19);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_33 = _zz_stateReg_17;
    end else begin
      _zz_stateReg_33 = (((_zz_stateReg_16 ^ (_zz_stateReg_17[7] ? (_zz_stateReg_62 ^ 8'h1b) : _zz_stateReg_62)) ^ ((_zz_stateReg_18[7] ? (_zz_stateReg_63 ^ 8'h1b) : _zz_stateReg_63) ^ _zz_stateReg_18)) ^ _zz_stateReg_19);
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_34 = _zz_stateReg_18;
    end else begin
      _zz_stateReg_34 = (((_zz_stateReg_16 ^ _zz_stateReg_17) ^ (_zz_stateReg_18[7] ? (_zz_stateReg_64 ^ 8'h1b) : _zz_stateReg_64)) ^ ((_zz_stateReg_19[7] ? (_zz_stateReg_65 ^ 8'h1b) : _zz_stateReg_65) ^ _zz_stateReg_19));
    end
  end

  always @(*) begin
    if(when_AES128_l272) begin
      _zz_stateReg_35 = _zz_stateReg_19;
    end else begin
      _zz_stateReg_35 = (((((_zz_stateReg_16[7] ? (_zz_stateReg_66 ^ 8'h1b) : _zz_stateReg_66) ^ _zz_stateReg_16) ^ _zz_stateReg_17) ^ _zz_stateReg_18) ^ (_zz_stateReg_19[7] ? (_zz_stateReg_67 ^ 8'h1b) : _zz_stateReg_67));
    end
  end

  assign _zz_stateReg_36 = _zz__zz_stateReg_36[7 : 0];
  assign _zz_stateReg_37 = _zz__zz_stateReg_37[7 : 0];
  assign _zz_stateReg_38 = _zz__zz_stateReg_38[7 : 0];
  assign _zz_stateReg_39 = _zz__zz_stateReg_39[7 : 0];
  assign _zz_stateReg_40 = _zz__zz_stateReg_40[7 : 0];
  assign _zz_stateReg_41 = _zz__zz_stateReg_41[7 : 0];
  assign _zz_stateReg_42 = _zz__zz_stateReg_42[7 : 0];
  assign _zz_stateReg_43 = _zz__zz_stateReg_43[7 : 0];
  assign _zz_stateReg_44 = _zz__zz_stateReg_44[7 : 0];
  assign _zz_stateReg_45 = _zz__zz_stateReg_45[7 : 0];
  assign _zz_stateReg_46 = _zz__zz_stateReg_46[7 : 0];
  assign _zz_stateReg_47 = _zz__zz_stateReg_47[7 : 0];
  assign _zz_stateReg_48 = _zz__zz_stateReg_48[7 : 0];
  assign _zz_stateReg_49 = _zz__zz_stateReg_49[7 : 0];
  assign _zz_stateReg_50 = _zz__zz_stateReg_50[7 : 0];
  assign _zz_stateReg_51 = _zz__zz_stateReg_51[7 : 0];
  assign _zz_stateReg_52 = _zz__zz_stateReg_52[7 : 0];
  assign _zz_stateReg_53 = _zz__zz_stateReg_53[7 : 0];
  assign _zz_stateReg_54 = _zz__zz_stateReg_54[7 : 0];
  assign _zz_stateReg_55 = _zz__zz_stateReg_55[7 : 0];
  assign _zz_stateReg_56 = _zz__zz_stateReg_56[7 : 0];
  assign _zz_stateReg_57 = _zz__zz_stateReg_57[7 : 0];
  assign _zz_stateReg_58 = _zz__zz_stateReg_58[7 : 0];
  assign _zz_stateReg_59 = _zz__zz_stateReg_59[7 : 0];
  assign _zz_stateReg_60 = _zz__zz_stateReg_60[7 : 0];
  assign _zz_stateReg_61 = _zz__zz_stateReg_61[7 : 0];
  assign _zz_stateReg_62 = _zz__zz_stateReg_62[7 : 0];
  assign _zz_stateReg_63 = _zz__zz_stateReg_63[7 : 0];
  assign _zz_stateReg_64 = _zz__zz_stateReg_64[7 : 0];
  assign _zz_stateReg_65 = _zz__zz_stateReg_65[7 : 0];
  assign _zz_stateReg_66 = _zz__zz_stateReg_66[7 : 0];
  assign _zz_stateReg_67 = _zz__zz_stateReg_67[7 : 0];
  assign _zz_stateReg_68 = {{{{{{{{{{{_zz__zz_stateReg_68,_zz__zz_stateReg_68_1},_zz_stateReg_26},_zz_stateReg_27},_zz_stateReg_28},_zz_stateReg_29},_zz_stateReg_30},_zz_stateReg_31},_zz_stateReg_32},_zz_stateReg_33},_zz_stateReg_34},_zz_stateReg_35};
  assign _zz_roundKeyReg_0 = _zz__zz_roundKeyReg_0;
  assign _zz_roundKeyReg_0_1 = {roundKeyReg_3[23 : 0],roundKeyReg_3[31 : 24]};
  assign _zz_roundKeyReg_0_2 = (roundKeyReg_0 ^ ({{{_zz__zz_roundKeyReg_0_2,_zz__zz_roundKeyReg_0_2_2},_zz__zz_roundKeyReg_0_2_4},_zz__zz_roundKeyReg_0_2_6} ^ {_zz_roundKeyReg_0,24'h0}));
  assign _zz_roundKeyReg_1 = (roundKeyReg_1 ^ _zz_roundKeyReg_0_2);
  assign _zz_roundKeyReg_2 = (roundKeyReg_2 ^ _zz_roundKeyReg_1);
  assign _zz_roundKeyReg_3 = (roundKeyReg_3 ^ _zz_roundKeyReg_2);
  assign _zz_stateReg_69 = {{{{{{{{{_zz__zz_stateReg_69,_zz__zz_stateReg_69_1},_zz__zz_stateReg_69_2},_zz_roundKeyReg_2[23 : 16]},_zz_roundKeyReg_2[15 : 8]},_zz_roundKeyReg_2[7 : 0]},_zz_roundKeyReg_3[31 : 24]},_zz_roundKeyReg_3[23 : 16]},_zz_roundKeyReg_3[15 : 8]},_zz_roundKeyReg_3[7 : 0]};
  assign when_AES128_l307 = (roundCount == 4'b1010);
  assign when_AES128_l313 = (rconCounter < 4'b1001);
  assign _zz_roundKeyReg_0_3 = io_key[127 : 96];
  assign _zz_roundKeyReg_1_1 = io_key[95 : 64];
  assign _zz_roundKeyReg_2_1 = io_key[63 : 32];
  assign _zz_roundKeyReg_3_1 = io_key[31 : 0];
  assign _zz_stateReg_70 = {roundKeyReg_3[23 : 0],roundKeyReg_3[31 : 24]};
  assign _zz_stateReg_71 = (roundKeyReg_0 ^ ({{{_zz__zz_stateReg_71,_zz__zz_stateReg_71_2},_zz__zz_stateReg_71_4},_zz__zz_stateReg_71_6} ^ {_zz__zz_stateReg_71_8,24'h0}));
  assign _zz_stateReg_72 = (roundKeyReg_1 ^ _zz_stateReg_71);
  assign _zz_stateReg_73 = (roundKeyReg_2 ^ _zz_stateReg_72);
  assign _zz_stateReg_74 = (roundKeyReg_3 ^ _zz_stateReg_73);
  assign when_AES128_l328 = (precomputeCounter == 4'b1001);
  assign _zz_roundKeyReg_3_2 = (roundKeyReg_3 ^ roundKeyReg_2);
  assign _zz_roundKeyReg_2_2 = (roundKeyReg_2 ^ roundKeyReg_1);
  assign _zz_roundKeyReg_1_2 = (roundKeyReg_1 ^ roundKeyReg_0);
  assign _zz_roundKeyReg_0_4 = {_zz_roundKeyReg_3_2[23 : 0],_zz_roundKeyReg_3_2[31 : 24]};
  assign _zz_roundKeyReg_0_5 = (roundKeyReg_0 ^ ({{{_zz__zz_roundKeyReg_0_5,_zz__zz_roundKeyReg_0_5_2},_zz__zz_roundKeyReg_0_5_4},_zz__zz_roundKeyReg_0_5_6} ^ {_zz_roundKeyReg_0,24'h0}));
  assign _zz_invMixed_0 = ({{{{{_zz__zz_invMixed_0,_zz__zz_invMixed_0_5},invSub_12},invSub_13},invSub_14},invSub_15} ^ {{{{{_zz__zz_invMixed_0_6,_zz__zz_invMixed_0_13},_zz__zz_invMixed_0_14},_zz_roundKeyReg_3_2[23 : 16]},_zz_roundKeyReg_3_2[15 : 8]},_zz_roundKeyReg_3_2[7 : 0]});
  assign _zz_invMixed_0_1 = _zz_invMixed_0[127 : 120];
  assign _zz_invMixed_0_2 = _zz_invMixed_0[119 : 112];
  assign _zz_invMixed_0_3 = _zz_invMixed_0[111 : 104];
  assign _zz_invMixed_0_4 = _zz_invMixed_0[103 : 96];
  assign _zz_invMixed_4 = _zz_invMixed_0[95 : 88];
  assign _zz_invMixed_4_1 = _zz_invMixed_0[87 : 80];
  assign _zz_invMixed_4_2 = _zz_invMixed_0[79 : 72];
  assign _zz_invMixed_4_3 = _zz_invMixed_0[71 : 64];
  assign _zz_invMixed_8 = _zz_invMixed_0[63 : 56];
  assign _zz_invMixed_8_1 = _zz_invMixed_0[55 : 48];
  assign _zz_invMixed_8_2 = _zz_invMixed_0[47 : 40];
  assign _zz_invMixed_8_3 = _zz_invMixed_0[39 : 32];
  assign _zz_invMixed_12 = _zz_invMixed_0[31 : 24];
  assign _zz_invMixed_12_1 = _zz_invMixed_0[23 : 16];
  assign _zz_invMixed_12_2 = _zz_invMixed_0[15 : 8];
  assign _zz_invMixed_12_3 = _zz_invMixed_0[7 : 0];
  assign when_AES128_l370 = (rconCounter == 4'b0000);
  assign _zz_invMixed_0_5 = _zz__zz_invMixed_0_5_1[7 : 0];
  assign _zz_invMixed_0_6 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_0_5 ^ 8'h1b) : _zz_invMixed_0_5);
  assign _zz_invMixed_0_7 = _zz__zz_invMixed_0_7_1[7 : 0];
  assign _zz_invMixed_0_8 = (_zz_invMixed_0_6[7] ? (_zz_invMixed_0_7 ^ 8'h1b) : _zz_invMixed_0_7);
  assign _zz_invMixed_0_9 = _zz__zz_invMixed_0_9_1[7 : 0];
  assign _zz_invMixed_0_10 = _zz__zz_invMixed_0_10_1[7 : 0];
  assign _zz_invMixed_0_11 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_0_10 ^ 8'h1b) : _zz_invMixed_0_10);
  assign _zz_invMixed_0_12 = _zz__zz_invMixed_0_12_1[7 : 0];
  assign _zz_invMixed_0_13 = _zz__zz_invMixed_0_13_1[7 : 0];
  assign _zz_invMixed_0_14 = _zz__zz_invMixed_0_14_1[7 : 0];
  assign _zz_invMixed_0_15 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_0_14 ^ 8'h1b) : _zz_invMixed_0_14);
  assign _zz_invMixed_0_16 = _zz__zz_invMixed_0_16[7 : 0];
  assign _zz_invMixed_0_17 = (_zz_invMixed_0_15[7] ? (_zz_invMixed_0_16 ^ 8'h1b) : _zz_invMixed_0_16);
  assign _zz_invMixed_0_18 = _zz__zz_invMixed_0_18[7 : 0];
  assign _zz_invMixed_0_19 = _zz__zz_invMixed_0_19[7 : 0];
  assign _zz_invMixed_0_20 = _zz__zz_invMixed_0_20[7 : 0];
  assign _zz_invMixed_0_21 = (_zz_invMixed_0_3[7] ? (_zz_invMixed_0_20 ^ 8'h1b) : _zz_invMixed_0_20);
  assign _zz_invMixed_0_22 = _zz__zz_invMixed_0_22[7 : 0];
  assign _zz_invMixed_0_23 = (_zz_invMixed_0_21[7] ? (_zz_invMixed_0_22 ^ 8'h1b) : _zz_invMixed_0_22);
  assign _zz_invMixed_0_24 = _zz__zz_invMixed_0_24[7 : 0];
  assign _zz_invMixed_0_25 = _zz__zz_invMixed_0_25[7 : 0];
  assign _zz_invMixed_0_26 = (_zz_invMixed_0_3[7] ? (_zz_invMixed_0_25 ^ 8'h1b) : _zz_invMixed_0_25);
  assign _zz_invMixed_0_27 = _zz__zz_invMixed_0_27[7 : 0];
  assign _zz_invMixed_0_28 = _zz__zz_invMixed_0_28[7 : 0];
  assign _zz_invMixed_0_29 = (_zz_invMixed_0_4[7] ? (_zz_invMixed_0_28 ^ 8'h1b) : _zz_invMixed_0_28);
  assign _zz_invMixed_0_30 = _zz__zz_invMixed_0_30[7 : 0];
  assign _zz_invMixed_0_31 = (_zz_invMixed_0_29[7] ? (_zz_invMixed_0_30 ^ 8'h1b) : _zz_invMixed_0_30);
  assign _zz_invMixed_0_32 = _zz__zz_invMixed_0_32[7 : 0];
  assign _zz_invMixed_1 = _zz__zz_invMixed_1[7 : 0];
  assign _zz_invMixed_1_1 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_1 ^ 8'h1b) : _zz_invMixed_1);
  assign _zz_invMixed_1_2 = _zz__zz_invMixed_1_2[7 : 0];
  assign _zz_invMixed_1_3 = (_zz_invMixed_1_1[7] ? (_zz_invMixed_1_2 ^ 8'h1b) : _zz_invMixed_1_2);
  assign _zz_invMixed_1_4 = _zz__zz_invMixed_1_4[7 : 0];
  assign _zz_invMixed_1_5 = _zz__zz_invMixed_1_5[7 : 0];
  assign _zz_invMixed_1_6 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_1_5 ^ 8'h1b) : _zz_invMixed_1_5);
  assign _zz_invMixed_1_7 = _zz__zz_invMixed_1_7[7 : 0];
  assign _zz_invMixed_1_8 = (_zz_invMixed_1_6[7] ? (_zz_invMixed_1_7 ^ 8'h1b) : _zz_invMixed_1_7);
  assign _zz_invMixed_1_9 = _zz__zz_invMixed_1_9[7 : 0];
  assign _zz_invMixed_1_10 = _zz__zz_invMixed_1_10[7 : 0];
  assign _zz_invMixed_1_11 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_1_10 ^ 8'h1b) : _zz_invMixed_1_10);
  assign _zz_invMixed_1_12 = _zz__zz_invMixed_1_12[7 : 0];
  assign _zz_invMixed_1_13 = _zz__zz_invMixed_1_13[7 : 0];
  assign _zz_invMixed_1_14 = _zz__zz_invMixed_1_14[7 : 0];
  assign _zz_invMixed_1_15 = (_zz_invMixed_0_3[7] ? (_zz_invMixed_1_14 ^ 8'h1b) : _zz_invMixed_1_14);
  assign _zz_invMixed_1_16 = _zz__zz_invMixed_1_16[7 : 0];
  assign _zz_invMixed_1_17 = (_zz_invMixed_1_15[7] ? (_zz_invMixed_1_16 ^ 8'h1b) : _zz_invMixed_1_16);
  assign _zz_invMixed_1_18 = _zz__zz_invMixed_1_18[7 : 0];
  assign _zz_invMixed_1_19 = _zz__zz_invMixed_1_19[7 : 0];
  assign _zz_invMixed_1_20 = _zz__zz_invMixed_1_20[7 : 0];
  assign _zz_invMixed_1_21 = (_zz_invMixed_0_4[7] ? (_zz_invMixed_1_20 ^ 8'h1b) : _zz_invMixed_1_20);
  assign _zz_invMixed_1_22 = _zz__zz_invMixed_1_22[7 : 0];
  assign _zz_invMixed_1_23 = (_zz_invMixed_1_21[7] ? (_zz_invMixed_1_22 ^ 8'h1b) : _zz_invMixed_1_22);
  assign _zz_invMixed_1_24 = _zz__zz_invMixed_1_24[7 : 0];
  assign _zz_invMixed_1_25 = _zz__zz_invMixed_1_25[7 : 0];
  assign _zz_invMixed_1_26 = (_zz_invMixed_0_4[7] ? (_zz_invMixed_1_25 ^ 8'h1b) : _zz_invMixed_1_25);
  assign _zz_invMixed_1_27 = _zz__zz_invMixed_1_27[7 : 0];
  assign _zz_invMixed_2 = _zz__zz_invMixed_2[7 : 0];
  assign _zz_invMixed_2_1 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_2 ^ 8'h1b) : _zz_invMixed_2);
  assign _zz_invMixed_2_2 = _zz__zz_invMixed_2_2[7 : 0];
  assign _zz_invMixed_2_3 = (_zz_invMixed_2_1[7] ? (_zz_invMixed_2_2 ^ 8'h1b) : _zz_invMixed_2_2);
  assign _zz_invMixed_2_4 = _zz__zz_invMixed_2_4[7 : 0];
  assign _zz_invMixed_2_5 = _zz__zz_invMixed_2_5[7 : 0];
  assign _zz_invMixed_2_6 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_2_5 ^ 8'h1b) : _zz_invMixed_2_5);
  assign _zz_invMixed_2_7 = _zz__zz_invMixed_2_7[7 : 0];
  assign _zz_invMixed_2_8 = _zz__zz_invMixed_2_8[7 : 0];
  assign _zz_invMixed_2_9 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_2_8 ^ 8'h1b) : _zz_invMixed_2_8);
  assign _zz_invMixed_2_10 = _zz__zz_invMixed_2_10[7 : 0];
  assign _zz_invMixed_2_11 = (_zz_invMixed_2_9[7] ? (_zz_invMixed_2_10 ^ 8'h1b) : _zz_invMixed_2_10);
  assign _zz_invMixed_2_12 = _zz__zz_invMixed_2_12[7 : 0];
  assign _zz_invMixed_2_13 = _zz__zz_invMixed_2_13[7 : 0];
  assign _zz_invMixed_2_14 = (_zz_invMixed_0_3[7] ? (_zz_invMixed_2_13 ^ 8'h1b) : _zz_invMixed_2_13);
  assign _zz_invMixed_2_15 = _zz__zz_invMixed_2_15[7 : 0];
  assign _zz_invMixed_2_16 = (_zz_invMixed_2_14[7] ? (_zz_invMixed_2_15 ^ 8'h1b) : _zz_invMixed_2_15);
  assign _zz_invMixed_2_17 = _zz__zz_invMixed_2_17[7 : 0];
  assign _zz_invMixed_2_18 = _zz__zz_invMixed_2_18[7 : 0];
  assign _zz_invMixed_2_19 = (_zz_invMixed_0_3[7] ? (_zz_invMixed_2_18 ^ 8'h1b) : _zz_invMixed_2_18);
  assign _zz_invMixed_2_20 = _zz__zz_invMixed_2_20[7 : 0];
  assign _zz_invMixed_2_21 = _zz__zz_invMixed_2_21[7 : 0];
  assign _zz_invMixed_2_22 = _zz__zz_invMixed_2_22[7 : 0];
  assign _zz_invMixed_2_23 = (_zz_invMixed_0_4[7] ? (_zz_invMixed_2_22 ^ 8'h1b) : _zz_invMixed_2_22);
  assign _zz_invMixed_2_24 = _zz__zz_invMixed_2_24[7 : 0];
  assign _zz_invMixed_2_25 = (_zz_invMixed_2_23[7] ? (_zz_invMixed_2_24 ^ 8'h1b) : _zz_invMixed_2_24);
  assign _zz_invMixed_2_26 = _zz__zz_invMixed_2_26[7 : 0];
  assign _zz_invMixed_2_27 = _zz__zz_invMixed_2_27[7 : 0];
  assign _zz_invMixed_3 = _zz__zz_invMixed_3[7 : 0];
  assign _zz_invMixed_3_1 = (_zz_invMixed_0_1[7] ? (_zz_invMixed_3 ^ 8'h1b) : _zz_invMixed_3);
  assign _zz_invMixed_3_2 = _zz__zz_invMixed_3_2[7 : 0];
  assign _zz_invMixed_3_3 = (_zz_invMixed_3_1[7] ? (_zz_invMixed_3_2 ^ 8'h1b) : _zz_invMixed_3_2);
  assign _zz_invMixed_3_4 = _zz__zz_invMixed_3_4[7 : 0];
  assign _zz_invMixed_3_5 = _zz__zz_invMixed_3_5[7 : 0];
  assign _zz_invMixed_3_6 = _zz__zz_invMixed_3_6[7 : 0];
  assign _zz_invMixed_3_7 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_3_6 ^ 8'h1b) : _zz_invMixed_3_6);
  assign _zz_invMixed_3_8 = _zz__zz_invMixed_3_8[7 : 0];
  assign _zz_invMixed_3_9 = (_zz_invMixed_3_7[7] ? (_zz_invMixed_3_8 ^ 8'h1b) : _zz_invMixed_3_8);
  assign _zz_invMixed_3_10 = _zz__zz_invMixed_3_10[7 : 0];
  assign _zz_invMixed_3_11 = _zz__zz_invMixed_3_11[7 : 0];
  assign _zz_invMixed_3_12 = (_zz_invMixed_0_2[7] ? (_zz_invMixed_3_11 ^ 8'h1b) : _zz_invMixed_3_11);
  assign _zz_invMixed_3_13 = _zz__zz_invMixed_3_13[7 : 0];
  assign _zz_invMixed_3_14 = _zz__zz_invMixed_3_14[7 : 0];
  assign _zz_invMixed_3_15 = (_zz_invMixed_0_3[7] ? (_zz_invMixed_3_14 ^ 8'h1b) : _zz_invMixed_3_14);
  assign _zz_invMixed_3_16 = _zz__zz_invMixed_3_16[7 : 0];
  assign _zz_invMixed_3_17 = (_zz_invMixed_3_15[7] ? (_zz_invMixed_3_16 ^ 8'h1b) : _zz_invMixed_3_16);
  assign _zz_invMixed_3_18 = _zz__zz_invMixed_3_18[7 : 0];
  assign _zz_invMixed_3_19 = _zz__zz_invMixed_3_19[7 : 0];
  assign _zz_invMixed_3_20 = (_zz_invMixed_0_4[7] ? (_zz_invMixed_3_19 ^ 8'h1b) : _zz_invMixed_3_19);
  assign _zz_invMixed_3_21 = _zz__zz_invMixed_3_21[7 : 0];
  assign _zz_invMixed_3_22 = (_zz_invMixed_3_20[7] ? (_zz_invMixed_3_21 ^ 8'h1b) : _zz_invMixed_3_21);
  assign _zz_invMixed_3_23 = _zz__zz_invMixed_3_23[7 : 0];
  assign _zz_invMixed_3_24 = _zz__zz_invMixed_3_24[7 : 0];
  assign _zz_invMixed_3_25 = (_zz_invMixed_0_4[7] ? (_zz_invMixed_3_24 ^ 8'h1b) : _zz_invMixed_3_24);
  assign _zz_invMixed_3_26 = _zz__zz_invMixed_3_26[7 : 0];
  assign _zz_invMixed_3_27 = _zz__zz_invMixed_3_27[7 : 0];
  assign _zz_invMixed_4_4 = _zz__zz_invMixed_4_4[7 : 0];
  assign _zz_invMixed_4_5 = (_zz_invMixed_4[7] ? (_zz_invMixed_4_4 ^ 8'h1b) : _zz_invMixed_4_4);
  assign _zz_invMixed_4_6 = _zz__zz_invMixed_4_6[7 : 0];
  assign _zz_invMixed_4_7 = (_zz_invMixed_4_5[7] ? (_zz_invMixed_4_6 ^ 8'h1b) : _zz_invMixed_4_6);
  assign _zz_invMixed_4_8 = _zz__zz_invMixed_4_8[7 : 0];
  assign _zz_invMixed_4_9 = _zz__zz_invMixed_4_9[7 : 0];
  assign _zz_invMixed_4_10 = (_zz_invMixed_4[7] ? (_zz_invMixed_4_9 ^ 8'h1b) : _zz_invMixed_4_9);
  assign _zz_invMixed_4_11 = _zz__zz_invMixed_4_11[7 : 0];
  assign _zz_invMixed_4_12 = _zz__zz_invMixed_4_12[7 : 0];
  assign _zz_invMixed_4_13 = _zz__zz_invMixed_4_13[7 : 0];
  assign _zz_invMixed_4_14 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_4_13 ^ 8'h1b) : _zz_invMixed_4_13);
  assign _zz_invMixed_4_15 = _zz__zz_invMixed_4_15[7 : 0];
  assign _zz_invMixed_4_16 = (_zz_invMixed_4_14[7] ? (_zz_invMixed_4_15 ^ 8'h1b) : _zz_invMixed_4_15);
  assign _zz_invMixed_4_17 = _zz__zz_invMixed_4_17[7 : 0];
  assign _zz_invMixed_4_18 = _zz__zz_invMixed_4_18[7 : 0];
  assign _zz_invMixed_4_19 = _zz__zz_invMixed_4_19[7 : 0];
  assign _zz_invMixed_4_20 = (_zz_invMixed_4_2[7] ? (_zz_invMixed_4_19 ^ 8'h1b) : _zz_invMixed_4_19);
  assign _zz_invMixed_4_21 = _zz__zz_invMixed_4_21[7 : 0];
  assign _zz_invMixed_4_22 = (_zz_invMixed_4_20[7] ? (_zz_invMixed_4_21 ^ 8'h1b) : _zz_invMixed_4_21);
  assign _zz_invMixed_4_23 = _zz__zz_invMixed_4_23[7 : 0];
  assign _zz_invMixed_4_24 = _zz__zz_invMixed_4_24[7 : 0];
  assign _zz_invMixed_4_25 = (_zz_invMixed_4_2[7] ? (_zz_invMixed_4_24 ^ 8'h1b) : _zz_invMixed_4_24);
  assign _zz_invMixed_4_26 = _zz__zz_invMixed_4_26[7 : 0];
  assign _zz_invMixed_4_27 = _zz__zz_invMixed_4_27[7 : 0];
  assign _zz_invMixed_4_28 = (_zz_invMixed_4_3[7] ? (_zz_invMixed_4_27 ^ 8'h1b) : _zz_invMixed_4_27);
  assign _zz_invMixed_4_29 = _zz__zz_invMixed_4_29[7 : 0];
  assign _zz_invMixed_4_30 = (_zz_invMixed_4_28[7] ? (_zz_invMixed_4_29 ^ 8'h1b) : _zz_invMixed_4_29);
  assign _zz_invMixed_4_31 = _zz__zz_invMixed_4_31[7 : 0];
  assign _zz_invMixed_5 = _zz__zz_invMixed_5[7 : 0];
  assign _zz_invMixed_5_1 = (_zz_invMixed_4[7] ? (_zz_invMixed_5 ^ 8'h1b) : _zz_invMixed_5);
  assign _zz_invMixed_5_2 = _zz__zz_invMixed_5_2[7 : 0];
  assign _zz_invMixed_5_3 = (_zz_invMixed_5_1[7] ? (_zz_invMixed_5_2 ^ 8'h1b) : _zz_invMixed_5_2);
  assign _zz_invMixed_5_4 = _zz__zz_invMixed_5_4[7 : 0];
  assign _zz_invMixed_5_5 = _zz__zz_invMixed_5_5[7 : 0];
  assign _zz_invMixed_5_6 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_5_5 ^ 8'h1b) : _zz_invMixed_5_5);
  assign _zz_invMixed_5_7 = _zz__zz_invMixed_5_7[7 : 0];
  assign _zz_invMixed_5_8 = (_zz_invMixed_5_6[7] ? (_zz_invMixed_5_7 ^ 8'h1b) : _zz_invMixed_5_7);
  assign _zz_invMixed_5_9 = _zz__zz_invMixed_5_9[7 : 0];
  assign _zz_invMixed_5_10 = _zz__zz_invMixed_5_10[7 : 0];
  assign _zz_invMixed_5_11 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_5_10 ^ 8'h1b) : _zz_invMixed_5_10);
  assign _zz_invMixed_5_12 = _zz__zz_invMixed_5_12[7 : 0];
  assign _zz_invMixed_5_13 = _zz__zz_invMixed_5_13[7 : 0];
  assign _zz_invMixed_5_14 = _zz__zz_invMixed_5_14[7 : 0];
  assign _zz_invMixed_5_15 = (_zz_invMixed_4_2[7] ? (_zz_invMixed_5_14 ^ 8'h1b) : _zz_invMixed_5_14);
  assign _zz_invMixed_5_16 = _zz__zz_invMixed_5_16[7 : 0];
  assign _zz_invMixed_5_17 = (_zz_invMixed_5_15[7] ? (_zz_invMixed_5_16 ^ 8'h1b) : _zz_invMixed_5_16);
  assign _zz_invMixed_5_18 = _zz__zz_invMixed_5_18[7 : 0];
  assign _zz_invMixed_5_19 = _zz__zz_invMixed_5_19[7 : 0];
  assign _zz_invMixed_5_20 = _zz__zz_invMixed_5_20[7 : 0];
  assign _zz_invMixed_5_21 = (_zz_invMixed_4_3[7] ? (_zz_invMixed_5_20 ^ 8'h1b) : _zz_invMixed_5_20);
  assign _zz_invMixed_5_22 = _zz__zz_invMixed_5_22[7 : 0];
  assign _zz_invMixed_5_23 = (_zz_invMixed_5_21[7] ? (_zz_invMixed_5_22 ^ 8'h1b) : _zz_invMixed_5_22);
  assign _zz_invMixed_5_24 = _zz__zz_invMixed_5_24[7 : 0];
  assign _zz_invMixed_5_25 = _zz__zz_invMixed_5_25[7 : 0];
  assign _zz_invMixed_5_26 = (_zz_invMixed_4_3[7] ? (_zz_invMixed_5_25 ^ 8'h1b) : _zz_invMixed_5_25);
  assign _zz_invMixed_5_27 = _zz__zz_invMixed_5_27[7 : 0];
  assign _zz_invMixed_6 = _zz__zz_invMixed_6[7 : 0];
  assign _zz_invMixed_6_1 = (_zz_invMixed_4[7] ? (_zz_invMixed_6 ^ 8'h1b) : _zz_invMixed_6);
  assign _zz_invMixed_6_2 = _zz__zz_invMixed_6_2[7 : 0];
  assign _zz_invMixed_6_3 = (_zz_invMixed_6_1[7] ? (_zz_invMixed_6_2 ^ 8'h1b) : _zz_invMixed_6_2);
  assign _zz_invMixed_6_4 = _zz__zz_invMixed_6_4[7 : 0];
  assign _zz_invMixed_6_5 = _zz__zz_invMixed_6_5[7 : 0];
  assign _zz_invMixed_6_6 = (_zz_invMixed_4[7] ? (_zz_invMixed_6_5 ^ 8'h1b) : _zz_invMixed_6_5);
  assign _zz_invMixed_6_7 = _zz__zz_invMixed_6_7[7 : 0];
  assign _zz_invMixed_6_8 = _zz__zz_invMixed_6_8[7 : 0];
  assign _zz_invMixed_6_9 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_6_8 ^ 8'h1b) : _zz_invMixed_6_8);
  assign _zz_invMixed_6_10 = _zz__zz_invMixed_6_10[7 : 0];
  assign _zz_invMixed_6_11 = (_zz_invMixed_6_9[7] ? (_zz_invMixed_6_10 ^ 8'h1b) : _zz_invMixed_6_10);
  assign _zz_invMixed_6_12 = _zz__zz_invMixed_6_12[7 : 0];
  assign _zz_invMixed_6_13 = _zz__zz_invMixed_6_13[7 : 0];
  assign _zz_invMixed_6_14 = (_zz_invMixed_4_2[7] ? (_zz_invMixed_6_13 ^ 8'h1b) : _zz_invMixed_6_13);
  assign _zz_invMixed_6_15 = _zz__zz_invMixed_6_15[7 : 0];
  assign _zz_invMixed_6_16 = (_zz_invMixed_6_14[7] ? (_zz_invMixed_6_15 ^ 8'h1b) : _zz_invMixed_6_15);
  assign _zz_invMixed_6_17 = _zz__zz_invMixed_6_17[7 : 0];
  assign _zz_invMixed_6_18 = _zz__zz_invMixed_6_18[7 : 0];
  assign _zz_invMixed_6_19 = (_zz_invMixed_4_2[7] ? (_zz_invMixed_6_18 ^ 8'h1b) : _zz_invMixed_6_18);
  assign _zz_invMixed_6_20 = _zz__zz_invMixed_6_20[7 : 0];
  assign _zz_invMixed_6_21 = _zz__zz_invMixed_6_21[7 : 0];
  assign _zz_invMixed_6_22 = _zz__zz_invMixed_6_22[7 : 0];
  assign _zz_invMixed_6_23 = (_zz_invMixed_4_3[7] ? (_zz_invMixed_6_22 ^ 8'h1b) : _zz_invMixed_6_22);
  assign _zz_invMixed_6_24 = _zz__zz_invMixed_6_24[7 : 0];
  assign _zz_invMixed_6_25 = (_zz_invMixed_6_23[7] ? (_zz_invMixed_6_24 ^ 8'h1b) : _zz_invMixed_6_24);
  assign _zz_invMixed_6_26 = _zz__zz_invMixed_6_26[7 : 0];
  assign _zz_invMixed_6_27 = _zz__zz_invMixed_6_27[7 : 0];
  assign _zz_invMixed_7 = _zz__zz_invMixed_7[7 : 0];
  assign _zz_invMixed_7_1 = (_zz_invMixed_4[7] ? (_zz_invMixed_7 ^ 8'h1b) : _zz_invMixed_7);
  assign _zz_invMixed_7_2 = _zz__zz_invMixed_7_2[7 : 0];
  assign _zz_invMixed_7_3 = (_zz_invMixed_7_1[7] ? (_zz_invMixed_7_2 ^ 8'h1b) : _zz_invMixed_7_2);
  assign _zz_invMixed_7_4 = _zz__zz_invMixed_7_4[7 : 0];
  assign _zz_invMixed_7_5 = _zz__zz_invMixed_7_5[7 : 0];
  assign _zz_invMixed_7_6 = _zz__zz_invMixed_7_6[7 : 0];
  assign _zz_invMixed_7_7 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_7_6 ^ 8'h1b) : _zz_invMixed_7_6);
  assign _zz_invMixed_7_8 = _zz__zz_invMixed_7_8[7 : 0];
  assign _zz_invMixed_7_9 = (_zz_invMixed_7_7[7] ? (_zz_invMixed_7_8 ^ 8'h1b) : _zz_invMixed_7_8);
  assign _zz_invMixed_7_10 = _zz__zz_invMixed_7_10[7 : 0];
  assign _zz_invMixed_7_11 = _zz__zz_invMixed_7_11[7 : 0];
  assign _zz_invMixed_7_12 = (_zz_invMixed_4_1[7] ? (_zz_invMixed_7_11 ^ 8'h1b) : _zz_invMixed_7_11);
  assign _zz_invMixed_7_13 = _zz__zz_invMixed_7_13[7 : 0];
  assign _zz_invMixed_7_14 = _zz__zz_invMixed_7_14[7 : 0];
  assign _zz_invMixed_7_15 = (_zz_invMixed_4_2[7] ? (_zz_invMixed_7_14 ^ 8'h1b) : _zz_invMixed_7_14);
  assign _zz_invMixed_7_16 = _zz__zz_invMixed_7_16[7 : 0];
  assign _zz_invMixed_7_17 = (_zz_invMixed_7_15[7] ? (_zz_invMixed_7_16 ^ 8'h1b) : _zz_invMixed_7_16);
  assign _zz_invMixed_7_18 = _zz__zz_invMixed_7_18[7 : 0];
  assign _zz_invMixed_7_19 = _zz__zz_invMixed_7_19[7 : 0];
  assign _zz_invMixed_7_20 = (_zz_invMixed_4_3[7] ? (_zz_invMixed_7_19 ^ 8'h1b) : _zz_invMixed_7_19);
  assign _zz_invMixed_7_21 = _zz__zz_invMixed_7_21[7 : 0];
  assign _zz_invMixed_7_22 = (_zz_invMixed_7_20[7] ? (_zz_invMixed_7_21 ^ 8'h1b) : _zz_invMixed_7_21);
  assign _zz_invMixed_7_23 = _zz__zz_invMixed_7_23[7 : 0];
  assign _zz_invMixed_7_24 = _zz__zz_invMixed_7_24[7 : 0];
  assign _zz_invMixed_7_25 = (_zz_invMixed_4_3[7] ? (_zz_invMixed_7_24 ^ 8'h1b) : _zz_invMixed_7_24);
  assign _zz_invMixed_7_26 = _zz__zz_invMixed_7_26[7 : 0];
  assign _zz_invMixed_7_27 = _zz__zz_invMixed_7_27[7 : 0];
  assign _zz_invMixed_8_4 = _zz__zz_invMixed_8_4[7 : 0];
  assign _zz_invMixed_8_5 = (_zz_invMixed_8[7] ? (_zz_invMixed_8_4 ^ 8'h1b) : _zz_invMixed_8_4);
  assign _zz_invMixed_8_6 = _zz__zz_invMixed_8_6[7 : 0];
  assign _zz_invMixed_8_7 = (_zz_invMixed_8_5[7] ? (_zz_invMixed_8_6 ^ 8'h1b) : _zz_invMixed_8_6);
  assign _zz_invMixed_8_8 = _zz__zz_invMixed_8_8[7 : 0];
  assign _zz_invMixed_8_9 = _zz__zz_invMixed_8_9[7 : 0];
  assign _zz_invMixed_8_10 = (_zz_invMixed_8[7] ? (_zz_invMixed_8_9 ^ 8'h1b) : _zz_invMixed_8_9);
  assign _zz_invMixed_8_11 = _zz__zz_invMixed_8_11[7 : 0];
  assign _zz_invMixed_8_12 = _zz__zz_invMixed_8_12[7 : 0];
  assign _zz_invMixed_8_13 = _zz__zz_invMixed_8_13[7 : 0];
  assign _zz_invMixed_8_14 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_8_13 ^ 8'h1b) : _zz_invMixed_8_13);
  assign _zz_invMixed_8_15 = _zz__zz_invMixed_8_15[7 : 0];
  assign _zz_invMixed_8_16 = (_zz_invMixed_8_14[7] ? (_zz_invMixed_8_15 ^ 8'h1b) : _zz_invMixed_8_15);
  assign _zz_invMixed_8_17 = _zz__zz_invMixed_8_17[7 : 0];
  assign _zz_invMixed_8_18 = _zz__zz_invMixed_8_18[7 : 0];
  assign _zz_invMixed_8_19 = _zz__zz_invMixed_8_19[7 : 0];
  assign _zz_invMixed_8_20 = (_zz_invMixed_8_2[7] ? (_zz_invMixed_8_19 ^ 8'h1b) : _zz_invMixed_8_19);
  assign _zz_invMixed_8_21 = _zz__zz_invMixed_8_21[7 : 0];
  assign _zz_invMixed_8_22 = (_zz_invMixed_8_20[7] ? (_zz_invMixed_8_21 ^ 8'h1b) : _zz_invMixed_8_21);
  assign _zz_invMixed_8_23 = _zz__zz_invMixed_8_23[7 : 0];
  assign _zz_invMixed_8_24 = _zz__zz_invMixed_8_24[7 : 0];
  assign _zz_invMixed_8_25 = (_zz_invMixed_8_2[7] ? (_zz_invMixed_8_24 ^ 8'h1b) : _zz_invMixed_8_24);
  assign _zz_invMixed_8_26 = _zz__zz_invMixed_8_26[7 : 0];
  assign _zz_invMixed_8_27 = _zz__zz_invMixed_8_27[7 : 0];
  assign _zz_invMixed_8_28 = (_zz_invMixed_8_3[7] ? (_zz_invMixed_8_27 ^ 8'h1b) : _zz_invMixed_8_27);
  assign _zz_invMixed_8_29 = _zz__zz_invMixed_8_29[7 : 0];
  assign _zz_invMixed_8_30 = (_zz_invMixed_8_28[7] ? (_zz_invMixed_8_29 ^ 8'h1b) : _zz_invMixed_8_29);
  assign _zz_invMixed_8_31 = _zz__zz_invMixed_8_31[7 : 0];
  assign _zz_invMixed_9 = _zz__zz_invMixed_9[7 : 0];
  assign _zz_invMixed_9_1 = (_zz_invMixed_8[7] ? (_zz_invMixed_9 ^ 8'h1b) : _zz_invMixed_9);
  assign _zz_invMixed_9_2 = _zz__zz_invMixed_9_2[7 : 0];
  assign _zz_invMixed_9_3 = (_zz_invMixed_9_1[7] ? (_zz_invMixed_9_2 ^ 8'h1b) : _zz_invMixed_9_2);
  assign _zz_invMixed_9_4 = _zz__zz_invMixed_9_4[7 : 0];
  assign _zz_invMixed_9_5 = _zz__zz_invMixed_9_5[7 : 0];
  assign _zz_invMixed_9_6 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_9_5 ^ 8'h1b) : _zz_invMixed_9_5);
  assign _zz_invMixed_9_7 = _zz__zz_invMixed_9_7[7 : 0];
  assign _zz_invMixed_9_8 = (_zz_invMixed_9_6[7] ? (_zz_invMixed_9_7 ^ 8'h1b) : _zz_invMixed_9_7);
  assign _zz_invMixed_9_9 = _zz__zz_invMixed_9_9[7 : 0];
  assign _zz_invMixed_9_10 = _zz__zz_invMixed_9_10[7 : 0];
  assign _zz_invMixed_9_11 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_9_10 ^ 8'h1b) : _zz_invMixed_9_10);
  assign _zz_invMixed_9_12 = _zz__zz_invMixed_9_12[7 : 0];
  assign _zz_invMixed_9_13 = _zz__zz_invMixed_9_13[7 : 0];
  assign _zz_invMixed_9_14 = _zz__zz_invMixed_9_14[7 : 0];
  assign _zz_invMixed_9_15 = (_zz_invMixed_8_2[7] ? (_zz_invMixed_9_14 ^ 8'h1b) : _zz_invMixed_9_14);
  assign _zz_invMixed_9_16 = _zz__zz_invMixed_9_16[7 : 0];
  assign _zz_invMixed_9_17 = (_zz_invMixed_9_15[7] ? (_zz_invMixed_9_16 ^ 8'h1b) : _zz_invMixed_9_16);
  assign _zz_invMixed_9_18 = _zz__zz_invMixed_9_18[7 : 0];
  assign _zz_invMixed_9_19 = _zz__zz_invMixed_9_19[7 : 0];
  assign _zz_invMixed_9_20 = _zz__zz_invMixed_9_20[7 : 0];
  assign _zz_invMixed_9_21 = (_zz_invMixed_8_3[7] ? (_zz_invMixed_9_20 ^ 8'h1b) : _zz_invMixed_9_20);
  assign _zz_invMixed_9_22 = _zz__zz_invMixed_9_22[7 : 0];
  assign _zz_invMixed_9_23 = (_zz_invMixed_9_21[7] ? (_zz_invMixed_9_22 ^ 8'h1b) : _zz_invMixed_9_22);
  assign _zz_invMixed_9_24 = _zz__zz_invMixed_9_24[7 : 0];
  assign _zz_invMixed_9_25 = _zz__zz_invMixed_9_25[7 : 0];
  assign _zz_invMixed_9_26 = (_zz_invMixed_8_3[7] ? (_zz_invMixed_9_25 ^ 8'h1b) : _zz_invMixed_9_25);
  assign _zz_invMixed_9_27 = _zz__zz_invMixed_9_27[7 : 0];
  assign _zz_invMixed_10 = _zz__zz_invMixed_10[7 : 0];
  assign _zz_invMixed_10_1 = (_zz_invMixed_8[7] ? (_zz_invMixed_10 ^ 8'h1b) : _zz_invMixed_10);
  assign _zz_invMixed_10_2 = _zz__zz_invMixed_10_2[7 : 0];
  assign _zz_invMixed_10_3 = (_zz_invMixed_10_1[7] ? (_zz_invMixed_10_2 ^ 8'h1b) : _zz_invMixed_10_2);
  assign _zz_invMixed_10_4 = _zz__zz_invMixed_10_4[7 : 0];
  assign _zz_invMixed_10_5 = _zz__zz_invMixed_10_5[7 : 0];
  assign _zz_invMixed_10_6 = (_zz_invMixed_8[7] ? (_zz_invMixed_10_5 ^ 8'h1b) : _zz_invMixed_10_5);
  assign _zz_invMixed_10_7 = _zz__zz_invMixed_10_7[7 : 0];
  assign _zz_invMixed_10_8 = _zz__zz_invMixed_10_8[7 : 0];
  assign _zz_invMixed_10_9 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_10_8 ^ 8'h1b) : _zz_invMixed_10_8);
  assign _zz_invMixed_10_10 = _zz__zz_invMixed_10_10[7 : 0];
  assign _zz_invMixed_10_11 = (_zz_invMixed_10_9[7] ? (_zz_invMixed_10_10 ^ 8'h1b) : _zz_invMixed_10_10);
  assign _zz_invMixed_10_12 = _zz__zz_invMixed_10_12[7 : 0];
  assign _zz_invMixed_10_13 = _zz__zz_invMixed_10_13[7 : 0];
  assign _zz_invMixed_10_14 = (_zz_invMixed_8_2[7] ? (_zz_invMixed_10_13 ^ 8'h1b) : _zz_invMixed_10_13);
  assign _zz_invMixed_10_15 = _zz__zz_invMixed_10_15[7 : 0];
  assign _zz_invMixed_10_16 = (_zz_invMixed_10_14[7] ? (_zz_invMixed_10_15 ^ 8'h1b) : _zz_invMixed_10_15);
  assign _zz_invMixed_10_17 = _zz__zz_invMixed_10_17[7 : 0];
  assign _zz_invMixed_10_18 = _zz__zz_invMixed_10_18[7 : 0];
  assign _zz_invMixed_10_19 = (_zz_invMixed_8_2[7] ? (_zz_invMixed_10_18 ^ 8'h1b) : _zz_invMixed_10_18);
  assign _zz_invMixed_10_20 = _zz__zz_invMixed_10_20[7 : 0];
  assign _zz_invMixed_10_21 = _zz__zz_invMixed_10_21[7 : 0];
  assign _zz_invMixed_10_22 = _zz__zz_invMixed_10_22[7 : 0];
  assign _zz_invMixed_10_23 = (_zz_invMixed_8_3[7] ? (_zz_invMixed_10_22 ^ 8'h1b) : _zz_invMixed_10_22);
  assign _zz_invMixed_10_24 = _zz__zz_invMixed_10_24[7 : 0];
  assign _zz_invMixed_10_25 = (_zz_invMixed_10_23[7] ? (_zz_invMixed_10_24 ^ 8'h1b) : _zz_invMixed_10_24);
  assign _zz_invMixed_10_26 = _zz__zz_invMixed_10_26[7 : 0];
  assign _zz_invMixed_10_27 = _zz__zz_invMixed_10_27[7 : 0];
  assign _zz_invMixed_11 = _zz__zz_invMixed_11[7 : 0];
  assign _zz_invMixed_11_1 = (_zz_invMixed_8[7] ? (_zz_invMixed_11 ^ 8'h1b) : _zz_invMixed_11);
  assign _zz_invMixed_11_2 = _zz__zz_invMixed_11_2[7 : 0];
  assign _zz_invMixed_11_3 = (_zz_invMixed_11_1[7] ? (_zz_invMixed_11_2 ^ 8'h1b) : _zz_invMixed_11_2);
  assign _zz_invMixed_11_4 = _zz__zz_invMixed_11_4[7 : 0];
  assign _zz_invMixed_11_5 = _zz__zz_invMixed_11_5[7 : 0];
  assign _zz_invMixed_11_6 = _zz__zz_invMixed_11_6[7 : 0];
  assign _zz_invMixed_11_7 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_11_6 ^ 8'h1b) : _zz_invMixed_11_6);
  assign _zz_invMixed_11_8 = _zz__zz_invMixed_11_8[7 : 0];
  assign _zz_invMixed_11_9 = (_zz_invMixed_11_7[7] ? (_zz_invMixed_11_8 ^ 8'h1b) : _zz_invMixed_11_8);
  assign _zz_invMixed_11_10 = _zz__zz_invMixed_11_10[7 : 0];
  assign _zz_invMixed_11_11 = _zz__zz_invMixed_11_11[7 : 0];
  assign _zz_invMixed_11_12 = (_zz_invMixed_8_1[7] ? (_zz_invMixed_11_11 ^ 8'h1b) : _zz_invMixed_11_11);
  assign _zz_invMixed_11_13 = _zz__zz_invMixed_11_13[7 : 0];
  assign _zz_invMixed_11_14 = _zz__zz_invMixed_11_14[7 : 0];
  assign _zz_invMixed_11_15 = (_zz_invMixed_8_2[7] ? (_zz_invMixed_11_14 ^ 8'h1b) : _zz_invMixed_11_14);
  assign _zz_invMixed_11_16 = _zz__zz_invMixed_11_16[7 : 0];
  assign _zz_invMixed_11_17 = (_zz_invMixed_11_15[7] ? (_zz_invMixed_11_16 ^ 8'h1b) : _zz_invMixed_11_16);
  assign _zz_invMixed_11_18 = _zz__zz_invMixed_11_18[7 : 0];
  assign _zz_invMixed_11_19 = _zz__zz_invMixed_11_19[7 : 0];
  assign _zz_invMixed_11_20 = (_zz_invMixed_8_3[7] ? (_zz_invMixed_11_19 ^ 8'h1b) : _zz_invMixed_11_19);
  assign _zz_invMixed_11_21 = _zz__zz_invMixed_11_21[7 : 0];
  assign _zz_invMixed_11_22 = (_zz_invMixed_11_20[7] ? (_zz_invMixed_11_21 ^ 8'h1b) : _zz_invMixed_11_21);
  assign _zz_invMixed_11_23 = _zz__zz_invMixed_11_23[7 : 0];
  assign _zz_invMixed_11_24 = _zz__zz_invMixed_11_24[7 : 0];
  assign _zz_invMixed_11_25 = (_zz_invMixed_8_3[7] ? (_zz_invMixed_11_24 ^ 8'h1b) : _zz_invMixed_11_24);
  assign _zz_invMixed_11_26 = _zz__zz_invMixed_11_26[7 : 0];
  assign _zz_invMixed_11_27 = _zz__zz_invMixed_11_27[7 : 0];
  assign _zz_invMixed_12_4 = _zz__zz_invMixed_12_4[7 : 0];
  assign _zz_invMixed_12_5 = (_zz_invMixed_12[7] ? (_zz_invMixed_12_4 ^ 8'h1b) : _zz_invMixed_12_4);
  assign _zz_invMixed_12_6 = _zz__zz_invMixed_12_6[7 : 0];
  assign _zz_invMixed_12_7 = (_zz_invMixed_12_5[7] ? (_zz_invMixed_12_6 ^ 8'h1b) : _zz_invMixed_12_6);
  assign _zz_invMixed_12_8 = _zz__zz_invMixed_12_8[7 : 0];
  assign _zz_invMixed_12_9 = _zz__zz_invMixed_12_9[7 : 0];
  assign _zz_invMixed_12_10 = (_zz_invMixed_12[7] ? (_zz_invMixed_12_9 ^ 8'h1b) : _zz_invMixed_12_9);
  assign _zz_invMixed_12_11 = _zz__zz_invMixed_12_11[7 : 0];
  assign _zz_invMixed_12_12 = _zz__zz_invMixed_12_12[7 : 0];
  assign _zz_invMixed_12_13 = _zz__zz_invMixed_12_13[7 : 0];
  assign _zz_invMixed_12_14 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_12_13 ^ 8'h1b) : _zz_invMixed_12_13);
  assign _zz_invMixed_12_15 = _zz__zz_invMixed_12_15[7 : 0];
  assign _zz_invMixed_12_16 = (_zz_invMixed_12_14[7] ? (_zz_invMixed_12_15 ^ 8'h1b) : _zz_invMixed_12_15);
  assign _zz_invMixed_12_17 = _zz__zz_invMixed_12_17[7 : 0];
  assign _zz_invMixed_12_18 = _zz__zz_invMixed_12_18[7 : 0];
  assign _zz_invMixed_12_19 = _zz__zz_invMixed_12_19[7 : 0];
  assign _zz_invMixed_12_20 = (_zz_invMixed_12_2[7] ? (_zz_invMixed_12_19 ^ 8'h1b) : _zz_invMixed_12_19);
  assign _zz_invMixed_12_21 = _zz__zz_invMixed_12_21[7 : 0];
  assign _zz_invMixed_12_22 = (_zz_invMixed_12_20[7] ? (_zz_invMixed_12_21 ^ 8'h1b) : _zz_invMixed_12_21);
  assign _zz_invMixed_12_23 = _zz__zz_invMixed_12_23[7 : 0];
  assign _zz_invMixed_12_24 = _zz__zz_invMixed_12_24[7 : 0];
  assign _zz_invMixed_12_25 = (_zz_invMixed_12_2[7] ? (_zz_invMixed_12_24 ^ 8'h1b) : _zz_invMixed_12_24);
  assign _zz_invMixed_12_26 = _zz__zz_invMixed_12_26[7 : 0];
  assign _zz_invMixed_12_27 = _zz__zz_invMixed_12_27[7 : 0];
  assign _zz_invMixed_12_28 = (_zz_invMixed_12_3[7] ? (_zz_invMixed_12_27 ^ 8'h1b) : _zz_invMixed_12_27);
  assign _zz_invMixed_12_29 = _zz__zz_invMixed_12_29[7 : 0];
  assign _zz_invMixed_12_30 = (_zz_invMixed_12_28[7] ? (_zz_invMixed_12_29 ^ 8'h1b) : _zz_invMixed_12_29);
  assign _zz_invMixed_12_31 = _zz__zz_invMixed_12_31[7 : 0];
  assign _zz_invMixed_13 = _zz__zz_invMixed_13[7 : 0];
  assign _zz_invMixed_13_1 = (_zz_invMixed_12[7] ? (_zz_invMixed_13 ^ 8'h1b) : _zz_invMixed_13);
  assign _zz_invMixed_13_2 = _zz__zz_invMixed_13_2[7 : 0];
  assign _zz_invMixed_13_3 = (_zz_invMixed_13_1[7] ? (_zz_invMixed_13_2 ^ 8'h1b) : _zz_invMixed_13_2);
  assign _zz_invMixed_13_4 = _zz__zz_invMixed_13_4[7 : 0];
  assign _zz_invMixed_13_5 = _zz__zz_invMixed_13_5[7 : 0];
  assign _zz_invMixed_13_6 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_13_5 ^ 8'h1b) : _zz_invMixed_13_5);
  assign _zz_invMixed_13_7 = _zz__zz_invMixed_13_7[7 : 0];
  assign _zz_invMixed_13_8 = (_zz_invMixed_13_6[7] ? (_zz_invMixed_13_7 ^ 8'h1b) : _zz_invMixed_13_7);
  assign _zz_invMixed_13_9 = _zz__zz_invMixed_13_9[7 : 0];
  assign _zz_invMixed_13_10 = _zz__zz_invMixed_13_10[7 : 0];
  assign _zz_invMixed_13_11 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_13_10 ^ 8'h1b) : _zz_invMixed_13_10);
  assign _zz_invMixed_13_12 = _zz__zz_invMixed_13_12[7 : 0];
  assign _zz_invMixed_13_13 = _zz__zz_invMixed_13_13[7 : 0];
  assign _zz_invMixed_13_14 = _zz__zz_invMixed_13_14[7 : 0];
  assign _zz_invMixed_13_15 = (_zz_invMixed_12_2[7] ? (_zz_invMixed_13_14 ^ 8'h1b) : _zz_invMixed_13_14);
  assign _zz_invMixed_13_16 = _zz__zz_invMixed_13_16[7 : 0];
  assign _zz_invMixed_13_17 = (_zz_invMixed_13_15[7] ? (_zz_invMixed_13_16 ^ 8'h1b) : _zz_invMixed_13_16);
  assign _zz_invMixed_13_18 = _zz__zz_invMixed_13_18[7 : 0];
  assign _zz_invMixed_13_19 = _zz__zz_invMixed_13_19[7 : 0];
  assign _zz_invMixed_13_20 = _zz__zz_invMixed_13_20[7 : 0];
  assign _zz_invMixed_13_21 = (_zz_invMixed_12_3[7] ? (_zz_invMixed_13_20 ^ 8'h1b) : _zz_invMixed_13_20);
  assign _zz_invMixed_13_22 = _zz__zz_invMixed_13_22[7 : 0];
  assign _zz_invMixed_13_23 = (_zz_invMixed_13_21[7] ? (_zz_invMixed_13_22 ^ 8'h1b) : _zz_invMixed_13_22);
  assign _zz_invMixed_13_24 = _zz__zz_invMixed_13_24[7 : 0];
  assign _zz_invMixed_13_25 = _zz__zz_invMixed_13_25[7 : 0];
  assign _zz_invMixed_13_26 = (_zz_invMixed_12_3[7] ? (_zz_invMixed_13_25 ^ 8'h1b) : _zz_invMixed_13_25);
  assign _zz_invMixed_13_27 = _zz__zz_invMixed_13_27[7 : 0];
  assign _zz_invMixed_14 = _zz__zz_invMixed_14[7 : 0];
  assign _zz_invMixed_14_1 = (_zz_invMixed_12[7] ? (_zz_invMixed_14 ^ 8'h1b) : _zz_invMixed_14);
  assign _zz_invMixed_14_2 = _zz__zz_invMixed_14_2[7 : 0];
  assign _zz_invMixed_14_3 = (_zz_invMixed_14_1[7] ? (_zz_invMixed_14_2 ^ 8'h1b) : _zz_invMixed_14_2);
  assign _zz_invMixed_14_4 = _zz__zz_invMixed_14_4[7 : 0];
  assign _zz_invMixed_14_5 = _zz__zz_invMixed_14_5[7 : 0];
  assign _zz_invMixed_14_6 = (_zz_invMixed_12[7] ? (_zz_invMixed_14_5 ^ 8'h1b) : _zz_invMixed_14_5);
  assign _zz_invMixed_14_7 = _zz__zz_invMixed_14_7[7 : 0];
  assign _zz_invMixed_14_8 = _zz__zz_invMixed_14_8[7 : 0];
  assign _zz_invMixed_14_9 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_14_8 ^ 8'h1b) : _zz_invMixed_14_8);
  assign _zz_invMixed_14_10 = _zz__zz_invMixed_14_10[7 : 0];
  assign _zz_invMixed_14_11 = (_zz_invMixed_14_9[7] ? (_zz_invMixed_14_10 ^ 8'h1b) : _zz_invMixed_14_10);
  assign _zz_invMixed_14_12 = _zz__zz_invMixed_14_12[7 : 0];
  assign _zz_invMixed_14_13 = _zz__zz_invMixed_14_13[7 : 0];
  assign _zz_invMixed_14_14 = (_zz_invMixed_12_2[7] ? (_zz_invMixed_14_13 ^ 8'h1b) : _zz_invMixed_14_13);
  assign _zz_invMixed_14_15 = _zz__zz_invMixed_14_15[7 : 0];
  assign _zz_invMixed_14_16 = (_zz_invMixed_14_14[7] ? (_zz_invMixed_14_15 ^ 8'h1b) : _zz_invMixed_14_15);
  assign _zz_invMixed_14_17 = _zz__zz_invMixed_14_17[7 : 0];
  assign _zz_invMixed_14_18 = _zz__zz_invMixed_14_18[7 : 0];
  assign _zz_invMixed_14_19 = (_zz_invMixed_12_2[7] ? (_zz_invMixed_14_18 ^ 8'h1b) : _zz_invMixed_14_18);
  assign _zz_invMixed_14_20 = _zz__zz_invMixed_14_20[7 : 0];
  assign _zz_invMixed_14_21 = _zz__zz_invMixed_14_21[7 : 0];
  assign _zz_invMixed_14_22 = _zz__zz_invMixed_14_22[7 : 0];
  assign _zz_invMixed_14_23 = (_zz_invMixed_12_3[7] ? (_zz_invMixed_14_22 ^ 8'h1b) : _zz_invMixed_14_22);
  assign _zz_invMixed_14_24 = _zz__zz_invMixed_14_24[7 : 0];
  assign _zz_invMixed_14_25 = (_zz_invMixed_14_23[7] ? (_zz_invMixed_14_24 ^ 8'h1b) : _zz_invMixed_14_24);
  assign _zz_invMixed_14_26 = _zz__zz_invMixed_14_26[7 : 0];
  assign _zz_invMixed_14_27 = _zz__zz_invMixed_14_27[7 : 0];
  assign _zz_invMixed_15 = _zz__zz_invMixed_15[7 : 0];
  assign _zz_invMixed_15_1 = (_zz_invMixed_12[7] ? (_zz_invMixed_15 ^ 8'h1b) : _zz_invMixed_15);
  assign _zz_invMixed_15_2 = _zz__zz_invMixed_15_2[7 : 0];
  assign _zz_invMixed_15_3 = (_zz_invMixed_15_1[7] ? (_zz_invMixed_15_2 ^ 8'h1b) : _zz_invMixed_15_2);
  assign _zz_invMixed_15_4 = _zz__zz_invMixed_15_4[7 : 0];
  assign _zz_invMixed_15_5 = _zz__zz_invMixed_15_5[7 : 0];
  assign _zz_invMixed_15_6 = _zz__zz_invMixed_15_6[7 : 0];
  assign _zz_invMixed_15_7 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_15_6 ^ 8'h1b) : _zz_invMixed_15_6);
  assign _zz_invMixed_15_8 = _zz__zz_invMixed_15_8[7 : 0];
  assign _zz_invMixed_15_9 = (_zz_invMixed_15_7[7] ? (_zz_invMixed_15_8 ^ 8'h1b) : _zz_invMixed_15_8);
  assign _zz_invMixed_15_10 = _zz__zz_invMixed_15_10[7 : 0];
  assign _zz_invMixed_15_11 = _zz__zz_invMixed_15_11[7 : 0];
  assign _zz_invMixed_15_12 = (_zz_invMixed_12_1[7] ? (_zz_invMixed_15_11 ^ 8'h1b) : _zz_invMixed_15_11);
  assign _zz_invMixed_15_13 = _zz__zz_invMixed_15_13[7 : 0];
  assign _zz_invMixed_15_14 = _zz__zz_invMixed_15_14[7 : 0];
  assign _zz_invMixed_15_15 = (_zz_invMixed_12_2[7] ? (_zz_invMixed_15_14 ^ 8'h1b) : _zz_invMixed_15_14);
  assign _zz_invMixed_15_16 = _zz__zz_invMixed_15_16[7 : 0];
  assign _zz_invMixed_15_17 = (_zz_invMixed_15_15[7] ? (_zz_invMixed_15_16 ^ 8'h1b) : _zz_invMixed_15_16);
  assign _zz_invMixed_15_18 = _zz__zz_invMixed_15_18[7 : 0];
  assign _zz_invMixed_15_19 = _zz__zz_invMixed_15_19[7 : 0];
  assign _zz_invMixed_15_20 = (_zz_invMixed_12_3[7] ? (_zz_invMixed_15_19 ^ 8'h1b) : _zz_invMixed_15_19);
  assign _zz_invMixed_15_21 = _zz__zz_invMixed_15_21[7 : 0];
  assign _zz_invMixed_15_22 = (_zz_invMixed_15_20[7] ? (_zz_invMixed_15_21 ^ 8'h1b) : _zz_invMixed_15_21);
  assign _zz_invMixed_15_23 = _zz__zz_invMixed_15_23[7 : 0];
  assign _zz_invMixed_15_24 = _zz__zz_invMixed_15_24[7 : 0];
  assign _zz_invMixed_15_25 = (_zz_invMixed_12_3[7] ? (_zz_invMixed_15_24 ^ 8'h1b) : _zz_invMixed_15_24);
  assign _zz_invMixed_15_26 = _zz__zz_invMixed_15_26[7 : 0];
  assign _zz_invMixed_15_27 = _zz__zz_invMixed_15_27[7 : 0];
  assign when_AES128_l397 = (roundCount == 4'b1010);
  assign when_AES128_l403 = (4'b0000 < rconCounter);
  assign when_AES128_l244 = (running && (! io_decrypt));
  assign when_AES128_l315 = (((! running) && (! precomputeRunning)) && io_decrypt);
  assign when_AES128_l339 = (running && io_decrypt);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      stateReg <= 128'h0;
      roundKeyReg_0 <= 32'h0;
      roundKeyReg_1 <= 32'h0;
      roundKeyReg_2 <= 32'h0;
      roundKeyReg_3 <= 32'h0;
      roundCount <= 4'b0000;
      running <= 1'b0;
      rconCounter <= 4'b0000;
      precomputeRunning <= 1'b0;
      precomputeCounter <= 4'b0000;
    end else begin
      if(when_AES128_l230) begin
        running <= 1'b1;
        stateReg <= {{{{{{_zz_stateReg_75,_zz_stateReg_87},_zz_stateReg_88},(_zz_stateReg_89 ^ _zz_stateReg_90)},(_zz_stateReg_91 ^ _zz_stateReg_3[23 : 16])},(io_dataIn[15 : 8] ^ _zz_stateReg_3[15 : 8])},(io_dataIn[7 : 0] ^ _zz_stateReg_3[7 : 0])};
        roundKeyReg_0 <= _zz_stateReg;
        roundKeyReg_1 <= _zz_stateReg_1;
        roundKeyReg_2 <= _zz_stateReg_2;
        roundKeyReg_3 <= _zz_stateReg_3;
        roundCount <= 4'b0000;
        rconCounter <= 4'b0000;
      end else begin
        if(when_AES128_l244) begin
          stateReg <= (_zz_stateReg_68 ^ _zz_stateReg_69);
          roundKeyReg_0 <= _zz_roundKeyReg_0_2;
          roundKeyReg_1 <= _zz_roundKeyReg_1;
          roundKeyReg_2 <= _zz_roundKeyReg_2;
          roundKeyReg_3 <= _zz_roundKeyReg_3;
          if(when_AES128_l307) begin
            running <= 1'b0;
          end else begin
            roundCount <= (roundCount + 4'b0001);
            if(when_AES128_l313) begin
              rconCounter <= (rconCounter + 4'b0001);
            end
          end
        end else begin
          if(when_AES128_l315) begin
            roundKeyReg_0 <= _zz_roundKeyReg_0_3;
            roundKeyReg_1 <= _zz_roundKeyReg_1_1;
            roundKeyReg_2 <= _zz_roundKeyReg_2_1;
            roundKeyReg_3 <= _zz_roundKeyReg_3_1;
            precomputeRunning <= 1'b1;
            precomputeCounter <= 4'b0000;
            rconCounter <= 4'b0000;
          end else begin
            if(precomputeRunning) begin
              roundKeyReg_0 <= _zz_stateReg_71;
              roundKeyReg_1 <= _zz_stateReg_72;
              roundKeyReg_2 <= _zz_stateReg_73;
              roundKeyReg_3 <= _zz_stateReg_74;
              precomputeCounter <= (precomputeCounter + 4'b0001);
              if(when_AES128_l328) begin
                precomputeRunning <= 1'b0;
                roundKeyReg_0 <= _zz_stateReg_71;
                roundKeyReg_1 <= _zz_stateReg_72;
                roundKeyReg_2 <= _zz_stateReg_73;
                roundKeyReg_3 <= _zz_stateReg_74;
                stateReg <= (io_dataIn ^ {{{{{{{{{_zz_stateReg_92,_zz_stateReg_93},_zz_stateReg_94},_zz_stateReg_73[23 : 16]},_zz_stateReg_73[15 : 8]},_zz_stateReg_73[7 : 0]},_zz_stateReg_74[31 : 24]},_zz_stateReg_74[23 : 16]},_zz_stateReg_74[15 : 8]},_zz_stateReg_74[7 : 0]});
                running <= 1'b1;
                roundCount <= 4'b0000;
                rconCounter <= 4'b1001;
              end
            end else begin
              if(when_AES128_l339) begin
                stateReg <= {{{{{{{{{{{_zz_stateReg_95,_zz_stateReg_96},invMixed_6},invMixed_7},invMixed_8},invMixed_9},invMixed_10},invMixed_11},invMixed_12},invMixed_13},invMixed_14},invMixed_15};
                roundKeyReg_0 <= _zz_roundKeyReg_0_5;
                roundKeyReg_1 <= _zz_roundKeyReg_1_2;
                roundKeyReg_2 <= _zz_roundKeyReg_2_2;
                roundKeyReg_3 <= _zz_roundKeyReg_3_2;
                if(when_AES128_l397) begin
                  running <= 1'b0;
                end else begin
                  roundCount <= (roundCount + 4'b0001);
                  if(when_AES128_l403) begin
                    rconCounter <= (rconCounter - 4'b0001);
                  end
                end
              end
            end
          end
        end
      end
    end
  end


endmodule
