// Generator : SpinalHDL v1.12.3    git head : 591e64062329e5e2e2b81f4d52422948053edb97
// Component : AesTop_WithAesIterative
// Git hash  : 1e0751b11cc7afb9e3f4716735fb6f9d1183579e

`timescale 1ns/1ps

module AesTop_WithAesIterative (
  input  wire          io_start,
  input  wire          io_decrypt,
  input  wire          io_key_bit,
  input  wire          io_dataIn_bit,
  output reg           io_dataOut_bit,
  output reg           io_busy,
  output reg           io_done,
  input  wire          io_clk,
  input  wire          io_reset
);

  reg                 area_aes_io_start;
  wire       [127:0]  area_aes_io_dataOut;
  wire                area_aes_io_busy;
  wire                area_aes_io_done;
  wire       [0:0]    _zz_area_keyExpanded;
  wire       [116:0]  _zz_area_keyExpanded_1;
  wire       [0:0]    _zz_area_keyExpanded_2;
  wire       [100:0]  _zz_area_keyExpanded_3;
  wire       [0:0]    _zz_area_keyExpanded_4;
  wire       [84:0]   _zz_area_keyExpanded_5;
  wire       [0:0]    _zz_area_keyExpanded_6;
  wire       [68:0]   _zz_area_keyExpanded_7;
  wire       [0:0]    _zz_area_keyExpanded_8;
  wire       [52:0]   _zz_area_keyExpanded_9;
  wire       [0:0]    _zz_area_keyExpanded_10;
  wire       [36:0]   _zz_area_keyExpanded_11;
  wire       [0:0]    _zz_area_keyExpanded_12;
  wire       [20:0]   _zz_area_keyExpanded_13;
  wire       [0:0]    _zz_area_keyExpanded_14;
  wire       [4:0]    _zz_area_keyExpanded_15;
  wire       [0:0]    _zz_area_dataExpanded;
  wire       [116:0]  _zz_area_dataExpanded_1;
  wire       [0:0]    _zz_area_dataExpanded_2;
  wire       [100:0]  _zz_area_dataExpanded_3;
  wire       [0:0]    _zz_area_dataExpanded_4;
  wire       [84:0]   _zz_area_dataExpanded_5;
  wire       [0:0]    _zz_area_dataExpanded_6;
  wire       [68:0]   _zz_area_dataExpanded_7;
  wire       [0:0]    _zz_area_dataExpanded_8;
  wire       [52:0]   _zz_area_dataExpanded_9;
  wire       [0:0]    _zz_area_dataExpanded_10;
  wire       [36:0]   _zz_area_dataExpanded_11;
  wire       [0:0]    _zz_area_dataExpanded_12;
  wire       [20:0]   _zz_area_dataExpanded_13;
  wire       [0:0]    _zz_area_dataExpanded_14;
  wire       [4:0]    _zz_area_dataExpanded_15;
  reg                 area_sampledKeyBit;
  reg                 area_sampledDataBit;
  wire       [127:0]  area_keyExpanded;
  wire       [127:0]  area_dataExpanded;
  reg        [1:0]    area_state;
  wire       [1:0]    area_IDLE;
  wire       [1:0]    area_START;
  wire       [1:0]    area_WAIT;
  wire       [1:0]    area_DONE;

  assign _zz_area_keyExpanded = area_sampledKeyBit;
  assign _zz_area_keyExpanded_1 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_2,_zz_area_keyExpanded_3}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_2 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_3 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_4,_zz_area_keyExpanded_5}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_4 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_5 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_6,_zz_area_keyExpanded_7}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_6 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_7 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_8,_zz_area_keyExpanded_9}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_8 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_9 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_10,_zz_area_keyExpanded_11}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_10 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_11 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_12,_zz_area_keyExpanded_13}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_12 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_13 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded_14,_zz_area_keyExpanded_15}}}}}}}}}}}}}}}};
  assign _zz_area_keyExpanded_14 = area_sampledKeyBit;
  assign _zz_area_keyExpanded_15 = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,area_sampledKeyBit}}}};
  assign _zz_area_dataExpanded = area_sampledDataBit;
  assign _zz_area_dataExpanded_1 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_2,_zz_area_dataExpanded_3}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_2 = area_sampledDataBit;
  assign _zz_area_dataExpanded_3 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_4,_zz_area_dataExpanded_5}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_4 = area_sampledDataBit;
  assign _zz_area_dataExpanded_5 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_6,_zz_area_dataExpanded_7}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_6 = area_sampledDataBit;
  assign _zz_area_dataExpanded_7 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_8,_zz_area_dataExpanded_9}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_8 = area_sampledDataBit;
  assign _zz_area_dataExpanded_9 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_10,_zz_area_dataExpanded_11}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_10 = area_sampledDataBit;
  assign _zz_area_dataExpanded_11 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_12,_zz_area_dataExpanded_13}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_12 = area_sampledDataBit;
  assign _zz_area_dataExpanded_13 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded_14,_zz_area_dataExpanded_15}}}}}}}}}}}}}}}};
  assign _zz_area_dataExpanded_14 = area_sampledDataBit;
  assign _zz_area_dataExpanded_15 = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,area_sampledDataBit}}}};
  AesIterative area_aes (
    .io_start   (area_aes_io_start         ), //i
    .io_decrypt (io_decrypt                ), //i
    .io_key     (area_keyExpanded[127:0]   ), //i
    .io_dataIn  (area_dataExpanded[127:0]  ), //i
    .io_dataOut (area_aes_io_dataOut[127:0]), //o
    .io_busy    (area_aes_io_busy          ), //o
    .io_done    (area_aes_io_done          ), //o
    .io_clk     (io_clk                    ), //i
    .io_reset   (io_reset                  )  //i
  );
  assign area_keyExpanded = {area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{area_sampledKeyBit,{_zz_area_keyExpanded,_zz_area_keyExpanded_1}}}}}}}}}}};
  assign area_dataExpanded = {area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{area_sampledDataBit,{_zz_area_dataExpanded,_zz_area_dataExpanded_1}}}}}}}}}}};
  assign area_IDLE = 2'b00;
  assign area_START = 2'b01;
  assign area_WAIT = 2'b10;
  assign area_DONE = 2'b11;
  always @(*) begin
    area_aes_io_start = 1'b0;
    if((area_state == area_IDLE)) begin
        if(io_start) begin
          area_aes_io_start = 1'b1;
        end
    end else if((area_state == area_START)) begin
    end else if((area_state == area_WAIT)) begin
    end else if((area_state == area_DONE)) begin
    end
  end

  always @(*) begin
    io_busy = 1'b0;
    if((area_state == area_IDLE)) begin
        if(io_start) begin
          io_busy = 1'b1;
        end
    end else if((area_state == area_START)) begin
        io_busy = 1'b1;
    end else if((area_state == area_WAIT)) begin
        io_busy = 1'b1;
    end else if((area_state == area_DONE)) begin
        io_busy = 1'b0;
    end
  end

  always @(*) begin
    io_done = 1'b0;
    if((area_state == area_IDLE)) begin
    end else if((area_state == area_START)) begin
    end else if((area_state == area_WAIT)) begin
    end else if((area_state == area_DONE)) begin
        io_done = 1'b1;
    end
  end

  always @(*) begin
    io_dataOut_bit = 1'b0;
    if((area_state == area_IDLE)) begin
    end else if((area_state == area_START)) begin
    end else if((area_state == area_WAIT)) begin
    end else if((area_state == area_DONE)) begin
        io_dataOut_bit = (^area_aes_io_dataOut);
    end
  end

  always @(posedge io_clk or posedge io_reset) begin
    if(io_reset) begin
      area_sampledKeyBit <= 1'b0;
      area_sampledDataBit <= 1'b0;
      area_state <= 2'b00;
    end else begin
      area_sampledKeyBit <= io_key_bit;
      area_sampledDataBit <= io_dataIn_bit;
      if((area_state == area_IDLE)) begin
          if(io_start) begin
            area_state <= area_START;
          end
      end else if((area_state == area_START)) begin
          area_state <= area_WAIT;
      end else if((area_state == area_WAIT)) begin
          if(area_aes_io_done) begin
            area_state <= area_DONE;
          end
      end else if((area_state == area_DONE)) begin
          area_state <= area_IDLE;
      end
    end
  end


endmodule

module AesIterative (
  input  wire          io_start,
  input  wire          io_decrypt,
  input  wire [127:0]  io_key,
  input  wire [127:0]  io_dataIn,
  output reg  [127:0]  io_dataOut,
  output wire          io_busy,
  output reg           io_done,
  input  wire          io_clk,
  input  wire          io_reset
);

  wire       [79:0]   _zz_stateReg_556;
  wire       [39:0]   _zz_stateReg_557;
  wire       [7:0]    _zz_stateReg_558;
  wire       [7:0]    _zz_stateReg_559;
  wire       [7:0]    _zz_stateReg_560;
  wire       [7:0]    _zz_stateReg_561;
  wire       [7:0]    _zz_stateReg_562;
  wire       [7:0]    _zz_stateReg_563;
  wire       [7:0]    _zz_stateReg_564;
  wire       [7:0]    _zz_stateReg_565;
  wire       [7:0]    _zz_stateReg_566;
  wire       [7:0]    _zz_stateReg_567;
  wire       [7:0]    _zz_stateReg_568;
  wire       [7:0]    _zz_stateReg_569;
  wire       [7:0]    _zz_stateReg_570;
  wire       [7:0]    _zz_stateReg_571;
  wire       [7:0]    _zz_stateReg_572;
  reg        [7:0]    _zz__zz_stateReg_4;
  wire       [7:0]    _zz__zz_stateReg_4_1;
  reg        [7:0]    _zz__zz_stateReg_8;
  wire       [7:0]    _zz__zz_stateReg_8_1;
  reg        [7:0]    _zz__zz_stateReg_12;
  wire       [7:0]    _zz__zz_stateReg_12_1;
  reg        [7:0]    _zz__zz_stateReg_16;
  wire       [7:0]    _zz__zz_stateReg_16_1;
  reg        [7:0]    _zz__zz_stateReg_5;
  wire       [7:0]    _zz__zz_stateReg_5_1;
  reg        [7:0]    _zz__zz_stateReg_9;
  wire       [7:0]    _zz__zz_stateReg_9_1;
  reg        [7:0]    _zz__zz_stateReg_13;
  wire       [7:0]    _zz__zz_stateReg_13_1;
  reg        [7:0]    _zz__zz_stateReg_17;
  wire       [7:0]    _zz__zz_stateReg_17_1;
  reg        [7:0]    _zz__zz_stateReg_6;
  wire       [7:0]    _zz__zz_stateReg_6_1;
  reg        [7:0]    _zz__zz_stateReg_10;
  wire       [7:0]    _zz__zz_stateReg_10_1;
  reg        [7:0]    _zz__zz_stateReg_14;
  wire       [7:0]    _zz__zz_stateReg_14_1;
  reg        [7:0]    _zz__zz_stateReg_18;
  wire       [7:0]    _zz__zz_stateReg_18_1;
  reg        [7:0]    _zz__zz_stateReg_7;
  wire       [7:0]    _zz__zz_stateReg_7_1;
  reg        [7:0]    _zz__zz_stateReg_11;
  wire       [7:0]    _zz__zz_stateReg_11_1;
  reg        [7:0]    _zz__zz_stateReg_15;
  wire       [7:0]    _zz__zz_stateReg_15_1;
  reg        [7:0]    _zz__zz_stateReg_19;
  wire       [7:0]    _zz__zz_stateReg_19_1;
  wire       [8:0]    _zz__zz_stateReg_36;
  wire       [8:0]    _zz__zz_stateReg_37;
  wire       [8:0]    _zz__zz_stateReg_38;
  wire       [8:0]    _zz__zz_stateReg_39;
  wire       [8:0]    _zz__zz_stateReg_40;
  wire       [8:0]    _zz__zz_stateReg_41;
  wire       [8:0]    _zz__zz_stateReg_42;
  wire       [8:0]    _zz__zz_stateReg_43;
  wire       [8:0]    _zz__zz_stateReg_44;
  wire       [8:0]    _zz__zz_stateReg_45;
  wire       [8:0]    _zz__zz_stateReg_46;
  wire       [8:0]    _zz__zz_stateReg_47;
  wire       [8:0]    _zz__zz_stateReg_48;
  wire       [8:0]    _zz__zz_stateReg_49;
  wire       [8:0]    _zz__zz_stateReg_50;
  wire       [8:0]    _zz__zz_stateReg_51;
  wire       [8:0]    _zz__zz_stateReg_52;
  wire       [8:0]    _zz__zz_stateReg_53;
  wire       [8:0]    _zz__zz_stateReg_54;
  wire       [8:0]    _zz__zz_stateReg_55;
  wire       [8:0]    _zz__zz_stateReg_56;
  wire       [8:0]    _zz__zz_stateReg_57;
  wire       [8:0]    _zz__zz_stateReg_58;
  wire       [8:0]    _zz__zz_stateReg_59;
  wire       [8:0]    _zz__zz_stateReg_60;
  wire       [8:0]    _zz__zz_stateReg_61;
  wire       [8:0]    _zz__zz_stateReg_62;
  wire       [8:0]    _zz__zz_stateReg_63;
  wire       [8:0]    _zz__zz_stateReg_64;
  wire       [8:0]    _zz__zz_stateReg_65;
  wire       [8:0]    _zz__zz_stateReg_66;
  wire       [8:0]    _zz__zz_stateReg_67;
  wire       [39:0]   _zz__zz_stateReg_68;
  wire       [7:0]    _zz__zz_stateReg_68_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_3;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2_4;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_5;
  reg        [7:0]    _zz__zz_roundKeyReg_0_2_6;
  wire       [7:0]    _zz__zz_roundKeyReg_0_2_7;
  wire       [55:0]   _zz__zz_stateReg_69;
  wire       [7:0]    _zz__zz_stateReg_69_1;
  wire       [7:0]    _zz__zz_stateReg_69_2;
  reg        [7:0]    _zz__zz_stateReg_71;
  wire       [7:0]    _zz__zz_stateReg_71_1;
  reg        [7:0]    _zz__zz_stateReg_71_2;
  wire       [7:0]    _zz__zz_stateReg_71_3;
  reg        [7:0]    _zz__zz_stateReg_71_4;
  wire       [7:0]    _zz__zz_stateReg_71_5;
  reg        [7:0]    _zz__zz_stateReg_71_6;
  wire       [7:0]    _zz__zz_stateReg_71_7;
  reg        [7:0]    _zz__zz_stateReg_71_8;
  wire       [55:0]   _zz_stateReg_573;
  wire       [7:0]    _zz_stateReg_574;
  wire       [7:0]    _zz_stateReg_575;
  reg        [7:0]    _zz__zz_roundKeyReg_0_4;
  wire       [7:0]    _zz__zz_roundKeyReg_0_4_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0_4_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_4_3;
  reg        [7:0]    _zz__zz_roundKeyReg_0_4_4;
  wire       [7:0]    _zz__zz_roundKeyReg_0_4_5;
  reg        [7:0]    _zz__zz_roundKeyReg_0_4_6;
  wire       [7:0]    _zz__zz_roundKeyReg_0_4_7;
  wire       [79:0]   _zz__zz_stateReg_75;
  wire       [31:0]   _zz__zz_stateReg_75_1;
  reg        [7:0]    _zz__zz_stateReg_75_2;
  wire       [7:0]    _zz__zz_stateReg_75_3;
  reg        [7:0]    _zz__zz_stateReg_75_4;
  wire       [7:0]    _zz__zz_stateReg_75_5;
  reg        [7:0]    _zz__zz_stateReg_75_6;
  wire       [7:0]    _zz__zz_stateReg_75_7;
  reg        [7:0]    _zz__zz_stateReg_75_8;
  wire       [7:0]    _zz__zz_stateReg_75_9;
  wire       [7:0]    _zz__zz_stateReg_75_10;
  reg        [7:0]    _zz__zz_stateReg_75_11;
  wire       [7:0]    _zz__zz_stateReg_75_12;
  reg        [7:0]    _zz__zz_stateReg_75_13;
  wire       [7:0]    _zz__zz_stateReg_75_14;
  reg        [7:0]    _zz__zz_stateReg_75_15;
  wire       [7:0]    _zz__zz_stateReg_75_16;
  reg        [7:0]    _zz__zz_stateReg_75_17;
  wire       [7:0]    _zz__zz_stateReg_75_18;
  reg        [7:0]    _zz__zz_stateReg_75_19;
  wire       [7:0]    _zz__zz_stateReg_75_20;
  reg        [7:0]    _zz__zz_stateReg_75_21;
  wire       [7:0]    _zz__zz_stateReg_75_22;
  wire       [7:0]    _zz__zz_stateReg_75_23;
  reg        [7:0]    _zz__zz_stateReg_75_24;
  wire       [7:0]    _zz__zz_stateReg_75_25;
  reg        [7:0]    _zz__zz_stateReg_75_26;
  wire       [7:0]    _zz__zz_stateReg_75_27;
  reg        [7:0]    _zz__zz_stateReg_75_28;
  wire       [7:0]    _zz__zz_stateReg_75_29;
  reg        [7:0]    _zz__zz_stateReg_75_30;
  wire       [7:0]    _zz__zz_stateReg_75_31;
  reg        [7:0]    _zz__zz_stateReg_75_32;
  wire       [7:0]    _zz__zz_stateReg_75_33;
  reg        [7:0]    _zz__zz_stateReg_75_34;
  wire       [7:0]    _zz__zz_stateReg_75_35;
  wire       [79:0]   _zz__zz_stateReg_75_36;
  wire       [31:0]   _zz__zz_stateReg_75_37;
  wire       [7:0]    _zz__zz_stateReg_75_38;
  wire       [7:0]    _zz__zz_stateReg_75_39;
  wire       [7:0]    _zz__zz_stateReg_75_40;
  wire       [7:0]    _zz__zz_stateReg_75_41;
  wire       [8:0]    _zz__zz_stateReg_108;
  wire       [8:0]    _zz__zz_stateReg_110;
  wire       [8:0]    _zz__zz_stateReg_112;
  wire       [8:0]    _zz__zz_stateReg_113;
  wire       [8:0]    _zz__zz_stateReg_115;
  wire       [8:0]    _zz__zz_stateReg_116;
  wire       [8:0]    _zz__zz_stateReg_117;
  wire       [8:0]    _zz__zz_stateReg_119;
  wire       [8:0]    _zz__zz_stateReg_121;
  wire       [8:0]    _zz__zz_stateReg_122;
  wire       [8:0]    _zz__zz_stateReg_123;
  wire       [8:0]    _zz__zz_stateReg_125;
  wire       [8:0]    _zz__zz_stateReg_127;
  wire       [8:0]    _zz__zz_stateReg_128;
  wire       [8:0]    _zz__zz_stateReg_130;
  wire       [8:0]    _zz__zz_stateReg_131;
  wire       [8:0]    _zz__zz_stateReg_133;
  wire       [8:0]    _zz__zz_stateReg_135;
  wire       [8:0]    _zz__zz_stateReg_136;
  wire       [8:0]    _zz__zz_stateReg_138;
  wire       [8:0]    _zz__zz_stateReg_140;
  wire       [8:0]    _zz__zz_stateReg_141;
  wire       [8:0]    _zz__zz_stateReg_143;
  wire       [8:0]    _zz__zz_stateReg_145;
  wire       [8:0]    _zz__zz_stateReg_146;
  wire       [8:0]    _zz__zz_stateReg_148;
  wire       [8:0]    _zz__zz_stateReg_149;
  wire       [8:0]    _zz__zz_stateReg_150;
  wire       [8:0]    _zz__zz_stateReg_152;
  wire       [8:0]    _zz__zz_stateReg_154;
  wire       [8:0]    _zz__zz_stateReg_155;
  wire       [8:0]    _zz__zz_stateReg_156;
  wire       [8:0]    _zz__zz_stateReg_158;
  wire       [8:0]    _zz__zz_stateReg_160;
  wire       [8:0]    _zz__zz_stateReg_161;
  wire       [8:0]    _zz__zz_stateReg_163;
  wire       [8:0]    _zz__zz_stateReg_164;
  wire       [8:0]    _zz__zz_stateReg_166;
  wire       [8:0]    _zz__zz_stateReg_168;
  wire       [8:0]    _zz__zz_stateReg_169;
  wire       [8:0]    _zz__zz_stateReg_171;
  wire       [8:0]    _zz__zz_stateReg_172;
  wire       [8:0]    _zz__zz_stateReg_174;
  wire       [8:0]    _zz__zz_stateReg_176;
  wire       [8:0]    _zz__zz_stateReg_177;
  wire       [8:0]    _zz__zz_stateReg_179;
  wire       [8:0]    _zz__zz_stateReg_181;
  wire       [8:0]    _zz__zz_stateReg_182;
  wire       [8:0]    _zz__zz_stateReg_184;
  wire       [8:0]    _zz__zz_stateReg_185;
  wire       [8:0]    _zz__zz_stateReg_186;
  wire       [8:0]    _zz__zz_stateReg_188;
  wire       [8:0]    _zz__zz_stateReg_190;
  wire       [8:0]    _zz__zz_stateReg_191;
  wire       [8:0]    _zz__zz_stateReg_192;
  wire       [8:0]    _zz__zz_stateReg_194;
  wire       [8:0]    _zz__zz_stateReg_196;
  wire       [8:0]    _zz__zz_stateReg_197;
  wire       [8:0]    _zz__zz_stateReg_198;
  wire       [8:0]    _zz__zz_stateReg_200;
  wire       [8:0]    _zz__zz_stateReg_202;
  wire       [8:0]    _zz__zz_stateReg_203;
  wire       [8:0]    _zz__zz_stateReg_205;
  wire       [8:0]    _zz__zz_stateReg_206;
  wire       [8:0]    _zz__zz_stateReg_208;
  wire       [8:0]    _zz__zz_stateReg_210;
  wire       [8:0]    _zz__zz_stateReg_211;
  wire       [8:0]    _zz__zz_stateReg_213;
  wire       [8:0]    _zz__zz_stateReg_215;
  wire       [8:0]    _zz__zz_stateReg_216;
  wire       [8:0]    _zz__zz_stateReg_218;
  wire       [8:0]    _zz__zz_stateReg_219;
  wire       [7:0]    _zz__zz_stateReg_92;
  wire       [7:0]    _zz__zz_stateReg_92_1;
  wire                _zz__zz_stateReg_92_2;
  wire       [7:0]    _zz__zz_stateReg_92_3;
  wire       [7:0]    _zz__zz_stateReg_92_4;
  wire       [7:0]    _zz__zz_stateReg_92_5;
  wire                _zz__zz_stateReg_92_6;
  wire       [7:0]    _zz__zz_stateReg_92_7;
  wire                _zz__zz_stateReg_92_8;
  wire       [7:0]    _zz__zz_stateReg_92_9;
  wire                _zz__zz_stateReg_93;
  wire       [7:0]    _zz__zz_stateReg_93_1;
  wire       [7:0]    _zz__zz_stateReg_93_2;
  wire       [7:0]    _zz__zz_stateReg_93_3;
  wire                _zz__zz_stateReg_93_4;
  wire       [7:0]    _zz__zz_stateReg_93_5;
  wire                _zz__zz_stateReg_93_6;
  wire       [7:0]    _zz__zz_stateReg_93_7;
  wire                _zz__zz_stateReg_93_8;
  wire       [7:0]    _zz__zz_stateReg_93_9;
  wire       [7:0]    _zz__zz_stateReg_93_10;
  wire       [7:0]    _zz__zz_stateReg_93_11;
  wire       [7:0]    _zz__zz_stateReg_94;
  wire       [7:0]    _zz__zz_stateReg_94_1;
  wire                _zz__zz_stateReg_94_2;
  wire       [7:0]    _zz__zz_stateReg_94_3;
  wire                _zz__zz_stateReg_94_4;
  wire       [7:0]    _zz__zz_stateReg_94_5;
  wire                _zz__zz_stateReg_94_6;
  wire       [7:0]    _zz__zz_stateReg_94_7;
  wire       [7:0]    _zz__zz_stateReg_94_8;
  wire       [7:0]    _zz__zz_stateReg_94_9;
  wire       [7:0]    _zz__zz_stateReg_94_10;
  wire       [7:0]    _zz__zz_stateReg_95;
  wire       [7:0]    _zz__zz_stateReg_95_1;
  wire       [7:0]    _zz__zz_stateReg_95_2;
  wire       [7:0]    _zz__zz_stateReg_95_3;
  wire       [7:0]    _zz__zz_stateReg_95_4;
  wire       [7:0]    _zz__zz_stateReg_95_5;
  wire       [7:0]    _zz__zz_stateReg_95_6;
  wire       [8:0]    _zz__zz_stateReg_220;
  wire       [8:0]    _zz__zz_stateReg_222;
  wire       [8:0]    _zz__zz_stateReg_224;
  wire       [8:0]    _zz__zz_stateReg_225;
  wire       [8:0]    _zz__zz_stateReg_227;
  wire       [8:0]    _zz__zz_stateReg_228;
  wire       [8:0]    _zz__zz_stateReg_229;
  wire       [8:0]    _zz__zz_stateReg_231;
  wire       [8:0]    _zz__zz_stateReg_233;
  wire       [8:0]    _zz__zz_stateReg_234;
  wire       [8:0]    _zz__zz_stateReg_235;
  wire       [8:0]    _zz__zz_stateReg_237;
  wire       [8:0]    _zz__zz_stateReg_239;
  wire       [8:0]    _zz__zz_stateReg_240;
  wire       [8:0]    _zz__zz_stateReg_242;
  wire       [8:0]    _zz__zz_stateReg_243;
  wire       [8:0]    _zz__zz_stateReg_245;
  wire       [8:0]    _zz__zz_stateReg_247;
  wire       [8:0]    _zz__zz_stateReg_248;
  wire       [8:0]    _zz__zz_stateReg_250;
  wire       [8:0]    _zz__zz_stateReg_252;
  wire       [8:0]    _zz__zz_stateReg_253;
  wire       [8:0]    _zz__zz_stateReg_255;
  wire       [8:0]    _zz__zz_stateReg_257;
  wire       [8:0]    _zz__zz_stateReg_258;
  wire       [8:0]    _zz__zz_stateReg_260;
  wire       [8:0]    _zz__zz_stateReg_261;
  wire       [8:0]    _zz__zz_stateReg_262;
  wire       [8:0]    _zz__zz_stateReg_264;
  wire       [8:0]    _zz__zz_stateReg_266;
  wire       [8:0]    _zz__zz_stateReg_267;
  wire       [8:0]    _zz__zz_stateReg_268;
  wire       [8:0]    _zz__zz_stateReg_270;
  wire       [8:0]    _zz__zz_stateReg_272;
  wire       [8:0]    _zz__zz_stateReg_273;
  wire       [8:0]    _zz__zz_stateReg_275;
  wire       [8:0]    _zz__zz_stateReg_276;
  wire       [8:0]    _zz__zz_stateReg_278;
  wire       [8:0]    _zz__zz_stateReg_280;
  wire       [8:0]    _zz__zz_stateReg_281;
  wire       [8:0]    _zz__zz_stateReg_283;
  wire       [8:0]    _zz__zz_stateReg_284;
  wire       [8:0]    _zz__zz_stateReg_286;
  wire       [8:0]    _zz__zz_stateReg_288;
  wire       [8:0]    _zz__zz_stateReg_289;
  wire       [8:0]    _zz__zz_stateReg_291;
  wire       [8:0]    _zz__zz_stateReg_293;
  wire       [8:0]    _zz__zz_stateReg_294;
  wire       [8:0]    _zz__zz_stateReg_296;
  wire       [8:0]    _zz__zz_stateReg_297;
  wire       [8:0]    _zz__zz_stateReg_298;
  wire       [8:0]    _zz__zz_stateReg_300;
  wire       [8:0]    _zz__zz_stateReg_302;
  wire       [8:0]    _zz__zz_stateReg_303;
  wire       [8:0]    _zz__zz_stateReg_304;
  wire       [8:0]    _zz__zz_stateReg_306;
  wire       [8:0]    _zz__zz_stateReg_308;
  wire       [8:0]    _zz__zz_stateReg_309;
  wire       [8:0]    _zz__zz_stateReg_310;
  wire       [8:0]    _zz__zz_stateReg_312;
  wire       [8:0]    _zz__zz_stateReg_314;
  wire       [8:0]    _zz__zz_stateReg_315;
  wire       [8:0]    _zz__zz_stateReg_317;
  wire       [8:0]    _zz__zz_stateReg_318;
  wire       [8:0]    _zz__zz_stateReg_320;
  wire       [8:0]    _zz__zz_stateReg_322;
  wire       [8:0]    _zz__zz_stateReg_323;
  wire       [8:0]    _zz__zz_stateReg_325;
  wire       [8:0]    _zz__zz_stateReg_327;
  wire       [8:0]    _zz__zz_stateReg_328;
  wire       [8:0]    _zz__zz_stateReg_330;
  wire       [8:0]    _zz__zz_stateReg_331;
  wire       [7:0]    _zz__zz_stateReg_96;
  wire       [7:0]    _zz__zz_stateReg_96_1;
  wire                _zz__zz_stateReg_96_2;
  wire       [7:0]    _zz__zz_stateReg_96_3;
  wire       [7:0]    _zz__zz_stateReg_96_4;
  wire       [7:0]    _zz__zz_stateReg_96_5;
  wire                _zz__zz_stateReg_96_6;
  wire       [7:0]    _zz__zz_stateReg_96_7;
  wire                _zz__zz_stateReg_96_8;
  wire       [7:0]    _zz__zz_stateReg_96_9;
  wire                _zz__zz_stateReg_97;
  wire       [7:0]    _zz__zz_stateReg_97_1;
  wire       [7:0]    _zz__zz_stateReg_97_2;
  wire       [7:0]    _zz__zz_stateReg_97_3;
  wire                _zz__zz_stateReg_97_4;
  wire       [7:0]    _zz__zz_stateReg_97_5;
  wire                _zz__zz_stateReg_97_6;
  wire       [7:0]    _zz__zz_stateReg_97_7;
  wire                _zz__zz_stateReg_97_8;
  wire       [7:0]    _zz__zz_stateReg_97_9;
  wire       [7:0]    _zz__zz_stateReg_97_10;
  wire       [7:0]    _zz__zz_stateReg_97_11;
  wire       [7:0]    _zz__zz_stateReg_98;
  wire       [7:0]    _zz__zz_stateReg_98_1;
  wire                _zz__zz_stateReg_98_2;
  wire       [7:0]    _zz__zz_stateReg_98_3;
  wire                _zz__zz_stateReg_98_4;
  wire       [7:0]    _zz__zz_stateReg_98_5;
  wire                _zz__zz_stateReg_98_6;
  wire       [7:0]    _zz__zz_stateReg_98_7;
  wire       [7:0]    _zz__zz_stateReg_98_8;
  wire       [7:0]    _zz__zz_stateReg_98_9;
  wire       [7:0]    _zz__zz_stateReg_98_10;
  wire       [7:0]    _zz__zz_stateReg_99;
  wire       [7:0]    _zz__zz_stateReg_99_1;
  wire       [7:0]    _zz__zz_stateReg_99_2;
  wire       [7:0]    _zz__zz_stateReg_99_3;
  wire       [7:0]    _zz__zz_stateReg_99_4;
  wire       [7:0]    _zz__zz_stateReg_99_5;
  wire       [7:0]    _zz__zz_stateReg_99_6;
  wire       [8:0]    _zz__zz_stateReg_332;
  wire       [8:0]    _zz__zz_stateReg_334;
  wire       [8:0]    _zz__zz_stateReg_336;
  wire       [8:0]    _zz__zz_stateReg_337;
  wire       [8:0]    _zz__zz_stateReg_339;
  wire       [8:0]    _zz__zz_stateReg_340;
  wire       [8:0]    _zz__zz_stateReg_341;
  wire       [8:0]    _zz__zz_stateReg_343;
  wire       [8:0]    _zz__zz_stateReg_345;
  wire       [8:0]    _zz__zz_stateReg_346;
  wire       [8:0]    _zz__zz_stateReg_347;
  wire       [8:0]    _zz__zz_stateReg_349;
  wire       [8:0]    _zz__zz_stateReg_351;
  wire       [8:0]    _zz__zz_stateReg_352;
  wire       [8:0]    _zz__zz_stateReg_354;
  wire       [8:0]    _zz__zz_stateReg_355;
  wire       [8:0]    _zz__zz_stateReg_357;
  wire       [8:0]    _zz__zz_stateReg_359;
  wire       [8:0]    _zz__zz_stateReg_360;
  wire       [8:0]    _zz__zz_stateReg_362;
  wire       [8:0]    _zz__zz_stateReg_364;
  wire       [8:0]    _zz__zz_stateReg_365;
  wire       [8:0]    _zz__zz_stateReg_367;
  wire       [8:0]    _zz__zz_stateReg_369;
  wire       [8:0]    _zz__zz_stateReg_370;
  wire       [8:0]    _zz__zz_stateReg_372;
  wire       [8:0]    _zz__zz_stateReg_373;
  wire       [8:0]    _zz__zz_stateReg_374;
  wire       [8:0]    _zz__zz_stateReg_376;
  wire       [8:0]    _zz__zz_stateReg_378;
  wire       [8:0]    _zz__zz_stateReg_379;
  wire       [8:0]    _zz__zz_stateReg_380;
  wire       [8:0]    _zz__zz_stateReg_382;
  wire       [8:0]    _zz__zz_stateReg_384;
  wire       [8:0]    _zz__zz_stateReg_385;
  wire       [8:0]    _zz__zz_stateReg_387;
  wire       [8:0]    _zz__zz_stateReg_388;
  wire       [8:0]    _zz__zz_stateReg_390;
  wire       [8:0]    _zz__zz_stateReg_392;
  wire       [8:0]    _zz__zz_stateReg_393;
  wire       [8:0]    _zz__zz_stateReg_395;
  wire       [8:0]    _zz__zz_stateReg_396;
  wire       [8:0]    _zz__zz_stateReg_398;
  wire       [8:0]    _zz__zz_stateReg_400;
  wire       [8:0]    _zz__zz_stateReg_401;
  wire       [8:0]    _zz__zz_stateReg_403;
  wire       [8:0]    _zz__zz_stateReg_405;
  wire       [8:0]    _zz__zz_stateReg_406;
  wire       [8:0]    _zz__zz_stateReg_408;
  wire       [8:0]    _zz__zz_stateReg_409;
  wire       [8:0]    _zz__zz_stateReg_410;
  wire       [8:0]    _zz__zz_stateReg_412;
  wire       [8:0]    _zz__zz_stateReg_414;
  wire       [8:0]    _zz__zz_stateReg_415;
  wire       [8:0]    _zz__zz_stateReg_416;
  wire       [8:0]    _zz__zz_stateReg_418;
  wire       [8:0]    _zz__zz_stateReg_420;
  wire       [8:0]    _zz__zz_stateReg_421;
  wire       [8:0]    _zz__zz_stateReg_422;
  wire       [8:0]    _zz__zz_stateReg_424;
  wire       [8:0]    _zz__zz_stateReg_426;
  wire       [8:0]    _zz__zz_stateReg_427;
  wire       [8:0]    _zz__zz_stateReg_429;
  wire       [8:0]    _zz__zz_stateReg_430;
  wire       [8:0]    _zz__zz_stateReg_432;
  wire       [8:0]    _zz__zz_stateReg_434;
  wire       [8:0]    _zz__zz_stateReg_435;
  wire       [8:0]    _zz__zz_stateReg_437;
  wire       [8:0]    _zz__zz_stateReg_439;
  wire       [8:0]    _zz__zz_stateReg_440;
  wire       [8:0]    _zz__zz_stateReg_442;
  wire       [8:0]    _zz__zz_stateReg_443;
  wire       [7:0]    _zz__zz_stateReg_100;
  wire       [7:0]    _zz__zz_stateReg_100_1;
  wire                _zz__zz_stateReg_100_2;
  wire       [7:0]    _zz__zz_stateReg_100_3;
  wire       [7:0]    _zz__zz_stateReg_100_4;
  wire       [7:0]    _zz__zz_stateReg_100_5;
  wire                _zz__zz_stateReg_100_6;
  wire       [7:0]    _zz__zz_stateReg_100_7;
  wire                _zz__zz_stateReg_100_8;
  wire       [7:0]    _zz__zz_stateReg_100_9;
  wire                _zz__zz_stateReg_101;
  wire       [7:0]    _zz__zz_stateReg_101_1;
  wire       [7:0]    _zz__zz_stateReg_101_2;
  wire       [7:0]    _zz__zz_stateReg_101_3;
  wire                _zz__zz_stateReg_101_4;
  wire       [7:0]    _zz__zz_stateReg_101_5;
  wire                _zz__zz_stateReg_101_6;
  wire       [7:0]    _zz__zz_stateReg_101_7;
  wire                _zz__zz_stateReg_101_8;
  wire       [7:0]    _zz__zz_stateReg_101_9;
  wire       [7:0]    _zz__zz_stateReg_101_10;
  wire       [7:0]    _zz__zz_stateReg_101_11;
  wire       [7:0]    _zz__zz_stateReg_102;
  wire       [7:0]    _zz__zz_stateReg_102_1;
  wire                _zz__zz_stateReg_102_2;
  wire       [7:0]    _zz__zz_stateReg_102_3;
  wire                _zz__zz_stateReg_102_4;
  wire       [7:0]    _zz__zz_stateReg_102_5;
  wire                _zz__zz_stateReg_102_6;
  wire       [7:0]    _zz__zz_stateReg_102_7;
  wire       [7:0]    _zz__zz_stateReg_102_8;
  wire       [7:0]    _zz__zz_stateReg_102_9;
  wire       [7:0]    _zz__zz_stateReg_102_10;
  wire       [7:0]    _zz__zz_stateReg_103;
  wire       [7:0]    _zz__zz_stateReg_103_1;
  wire       [7:0]    _zz__zz_stateReg_103_2;
  wire       [7:0]    _zz__zz_stateReg_103_3;
  wire       [7:0]    _zz__zz_stateReg_103_4;
  wire       [7:0]    _zz__zz_stateReg_103_5;
  wire       [7:0]    _zz__zz_stateReg_103_6;
  wire       [8:0]    _zz__zz_stateReg_444;
  wire       [8:0]    _zz__zz_stateReg_446;
  wire       [8:0]    _zz__zz_stateReg_448;
  wire       [8:0]    _zz__zz_stateReg_449;
  wire       [8:0]    _zz__zz_stateReg_451;
  wire       [8:0]    _zz__zz_stateReg_452;
  wire       [8:0]    _zz__zz_stateReg_453;
  wire       [8:0]    _zz__zz_stateReg_455;
  wire       [8:0]    _zz__zz_stateReg_457;
  wire       [8:0]    _zz__zz_stateReg_458;
  wire       [8:0]    _zz__zz_stateReg_459;
  wire       [8:0]    _zz__zz_stateReg_461;
  wire       [8:0]    _zz__zz_stateReg_463;
  wire       [8:0]    _zz__zz_stateReg_464;
  wire       [8:0]    _zz__zz_stateReg_466;
  wire       [8:0]    _zz__zz_stateReg_467;
  wire       [8:0]    _zz__zz_stateReg_469;
  wire       [8:0]    _zz__zz_stateReg_471;
  wire       [8:0]    _zz__zz_stateReg_472;
  wire       [8:0]    _zz__zz_stateReg_474;
  wire       [8:0]    _zz__zz_stateReg_476;
  wire       [8:0]    _zz__zz_stateReg_477;
  wire       [8:0]    _zz__zz_stateReg_479;
  wire       [8:0]    _zz__zz_stateReg_481;
  wire       [8:0]    _zz__zz_stateReg_482;
  wire       [8:0]    _zz__zz_stateReg_484;
  wire       [8:0]    _zz__zz_stateReg_485;
  wire       [8:0]    _zz__zz_stateReg_486;
  wire       [8:0]    _zz__zz_stateReg_488;
  wire       [8:0]    _zz__zz_stateReg_490;
  wire       [8:0]    _zz__zz_stateReg_491;
  wire       [8:0]    _zz__zz_stateReg_492;
  wire       [8:0]    _zz__zz_stateReg_494;
  wire       [8:0]    _zz__zz_stateReg_496;
  wire       [8:0]    _zz__zz_stateReg_497;
  wire       [8:0]    _zz__zz_stateReg_499;
  wire       [8:0]    _zz__zz_stateReg_500;
  wire       [8:0]    _zz__zz_stateReg_502;
  wire       [8:0]    _zz__zz_stateReg_504;
  wire       [8:0]    _zz__zz_stateReg_505;
  wire       [8:0]    _zz__zz_stateReg_507;
  wire       [8:0]    _zz__zz_stateReg_508;
  wire       [8:0]    _zz__zz_stateReg_510;
  wire       [8:0]    _zz__zz_stateReg_512;
  wire       [8:0]    _zz__zz_stateReg_513;
  wire       [8:0]    _zz__zz_stateReg_515;
  wire       [8:0]    _zz__zz_stateReg_517;
  wire       [8:0]    _zz__zz_stateReg_518;
  wire       [8:0]    _zz__zz_stateReg_520;
  wire       [8:0]    _zz__zz_stateReg_521;
  wire       [8:0]    _zz__zz_stateReg_522;
  wire       [8:0]    _zz__zz_stateReg_524;
  wire       [8:0]    _zz__zz_stateReg_526;
  wire       [8:0]    _zz__zz_stateReg_527;
  wire       [8:0]    _zz__zz_stateReg_528;
  wire       [8:0]    _zz__zz_stateReg_530;
  wire       [8:0]    _zz__zz_stateReg_532;
  wire       [8:0]    _zz__zz_stateReg_533;
  wire       [8:0]    _zz__zz_stateReg_534;
  wire       [8:0]    _zz__zz_stateReg_536;
  wire       [8:0]    _zz__zz_stateReg_538;
  wire       [8:0]    _zz__zz_stateReg_539;
  wire       [8:0]    _zz__zz_stateReg_541;
  wire       [8:0]    _zz__zz_stateReg_542;
  wire       [8:0]    _zz__zz_stateReg_544;
  wire       [8:0]    _zz__zz_stateReg_546;
  wire       [8:0]    _zz__zz_stateReg_547;
  wire       [8:0]    _zz__zz_stateReg_549;
  wire       [8:0]    _zz__zz_stateReg_551;
  wire       [8:0]    _zz__zz_stateReg_552;
  wire       [8:0]    _zz__zz_stateReg_554;
  wire       [8:0]    _zz__zz_stateReg_555;
  wire       [7:0]    _zz__zz_stateReg_104;
  wire       [7:0]    _zz__zz_stateReg_104_1;
  wire                _zz__zz_stateReg_104_2;
  wire       [7:0]    _zz__zz_stateReg_104_3;
  wire       [7:0]    _zz__zz_stateReg_104_4;
  wire       [7:0]    _zz__zz_stateReg_104_5;
  wire                _zz__zz_stateReg_104_6;
  wire       [7:0]    _zz__zz_stateReg_104_7;
  wire                _zz__zz_stateReg_104_8;
  wire       [7:0]    _zz__zz_stateReg_104_9;
  wire                _zz__zz_stateReg_105;
  wire       [7:0]    _zz__zz_stateReg_105_1;
  wire       [7:0]    _zz__zz_stateReg_105_2;
  wire       [7:0]    _zz__zz_stateReg_105_3;
  wire                _zz__zz_stateReg_105_4;
  wire       [7:0]    _zz__zz_stateReg_105_5;
  wire                _zz__zz_stateReg_105_6;
  wire       [7:0]    _zz__zz_stateReg_105_7;
  wire                _zz__zz_stateReg_105_8;
  wire       [7:0]    _zz__zz_stateReg_105_9;
  wire       [7:0]    _zz__zz_stateReg_105_10;
  wire       [7:0]    _zz__zz_stateReg_105_11;
  wire       [7:0]    _zz__zz_stateReg_106;
  wire       [7:0]    _zz__zz_stateReg_106_1;
  wire                _zz__zz_stateReg_106_2;
  wire       [7:0]    _zz__zz_stateReg_106_3;
  wire                _zz__zz_stateReg_106_4;
  wire       [7:0]    _zz__zz_stateReg_106_5;
  wire                _zz__zz_stateReg_106_6;
  wire       [7:0]    _zz__zz_stateReg_106_7;
  wire       [7:0]    _zz__zz_stateReg_106_8;
  wire       [7:0]    _zz__zz_stateReg_106_9;
  wire       [7:0]    _zz__zz_stateReg_106_10;
  wire       [7:0]    _zz__zz_stateReg_107;
  wire       [7:0]    _zz__zz_stateReg_107_1;
  wire       [7:0]    _zz__zz_stateReg_107_2;
  wire       [7:0]    _zz__zz_stateReg_107_3;
  wire       [7:0]    _zz__zz_stateReg_107_4;
  wire       [7:0]    _zz__zz_stateReg_107_5;
  wire       [7:0]    _zz__zz_stateReg_107_6;
  wire       [39:0]   _zz_stateReg_576;
  wire       [7:0]    _zz_stateReg_577;
  wire       [7:0]    rcon_0;
  wire       [7:0]    rcon_1;
  wire       [7:0]    rcon_2;
  wire       [7:0]    rcon_3;
  wire       [7:0]    rcon_4;
  wire       [7:0]    rcon_5;
  wire       [7:0]    rcon_6;
  wire       [7:0]    rcon_7;
  wire       [7:0]    rcon_8;
  wire       [7:0]    rcon_9;
  wire       [7:0]    sboxRom_0;
  wire       [7:0]    sboxRom_1;
  wire       [7:0]    sboxRom_2;
  wire       [7:0]    sboxRom_3;
  wire       [7:0]    sboxRom_4;
  wire       [7:0]    sboxRom_5;
  wire       [7:0]    sboxRom_6;
  wire       [7:0]    sboxRom_7;
  wire       [7:0]    sboxRom_8;
  wire       [7:0]    sboxRom_9;
  wire       [7:0]    sboxRom_10;
  wire       [7:0]    sboxRom_11;
  wire       [7:0]    sboxRom_12;
  wire       [7:0]    sboxRom_13;
  wire       [7:0]    sboxRom_14;
  wire       [7:0]    sboxRom_15;
  wire       [7:0]    sboxRom_16;
  wire       [7:0]    sboxRom_17;
  wire       [7:0]    sboxRom_18;
  wire       [7:0]    sboxRom_19;
  wire       [7:0]    sboxRom_20;
  wire       [7:0]    sboxRom_21;
  wire       [7:0]    sboxRom_22;
  wire       [7:0]    sboxRom_23;
  wire       [7:0]    sboxRom_24;
  wire       [7:0]    sboxRom_25;
  wire       [7:0]    sboxRom_26;
  wire       [7:0]    sboxRom_27;
  wire       [7:0]    sboxRom_28;
  wire       [7:0]    sboxRom_29;
  wire       [7:0]    sboxRom_30;
  wire       [7:0]    sboxRom_31;
  wire       [7:0]    sboxRom_32;
  wire       [7:0]    sboxRom_33;
  wire       [7:0]    sboxRom_34;
  wire       [7:0]    sboxRom_35;
  wire       [7:0]    sboxRom_36;
  wire       [7:0]    sboxRom_37;
  wire       [7:0]    sboxRom_38;
  wire       [7:0]    sboxRom_39;
  wire       [7:0]    sboxRom_40;
  wire       [7:0]    sboxRom_41;
  wire       [7:0]    sboxRom_42;
  wire       [7:0]    sboxRom_43;
  wire       [7:0]    sboxRom_44;
  wire       [7:0]    sboxRom_45;
  wire       [7:0]    sboxRom_46;
  wire       [7:0]    sboxRom_47;
  wire       [7:0]    sboxRom_48;
  wire       [7:0]    sboxRom_49;
  wire       [7:0]    sboxRom_50;
  wire       [7:0]    sboxRom_51;
  wire       [7:0]    sboxRom_52;
  wire       [7:0]    sboxRom_53;
  wire       [7:0]    sboxRom_54;
  wire       [7:0]    sboxRom_55;
  wire       [7:0]    sboxRom_56;
  wire       [7:0]    sboxRom_57;
  wire       [7:0]    sboxRom_58;
  wire       [7:0]    sboxRom_59;
  wire       [7:0]    sboxRom_60;
  wire       [7:0]    sboxRom_61;
  wire       [7:0]    sboxRom_62;
  wire       [7:0]    sboxRom_63;
  wire       [7:0]    sboxRom_64;
  wire       [7:0]    sboxRom_65;
  wire       [7:0]    sboxRom_66;
  wire       [7:0]    sboxRom_67;
  wire       [7:0]    sboxRom_68;
  wire       [7:0]    sboxRom_69;
  wire       [7:0]    sboxRom_70;
  wire       [7:0]    sboxRom_71;
  wire       [7:0]    sboxRom_72;
  wire       [7:0]    sboxRom_73;
  wire       [7:0]    sboxRom_74;
  wire       [7:0]    sboxRom_75;
  wire       [7:0]    sboxRom_76;
  wire       [7:0]    sboxRom_77;
  wire       [7:0]    sboxRom_78;
  wire       [7:0]    sboxRom_79;
  wire       [7:0]    sboxRom_80;
  wire       [7:0]    sboxRom_81;
  wire       [7:0]    sboxRom_82;
  wire       [7:0]    sboxRom_83;
  wire       [7:0]    sboxRom_84;
  wire       [7:0]    sboxRom_85;
  wire       [7:0]    sboxRom_86;
  wire       [7:0]    sboxRom_87;
  wire       [7:0]    sboxRom_88;
  wire       [7:0]    sboxRom_89;
  wire       [7:0]    sboxRom_90;
  wire       [7:0]    sboxRom_91;
  wire       [7:0]    sboxRom_92;
  wire       [7:0]    sboxRom_93;
  wire       [7:0]    sboxRom_94;
  wire       [7:0]    sboxRom_95;
  wire       [7:0]    sboxRom_96;
  wire       [7:0]    sboxRom_97;
  wire       [7:0]    sboxRom_98;
  wire       [7:0]    sboxRom_99;
  wire       [7:0]    sboxRom_100;
  wire       [7:0]    sboxRom_101;
  wire       [7:0]    sboxRom_102;
  wire       [7:0]    sboxRom_103;
  wire       [7:0]    sboxRom_104;
  wire       [7:0]    sboxRom_105;
  wire       [7:0]    sboxRom_106;
  wire       [7:0]    sboxRom_107;
  wire       [7:0]    sboxRom_108;
  wire       [7:0]    sboxRom_109;
  wire       [7:0]    sboxRom_110;
  wire       [7:0]    sboxRom_111;
  wire       [7:0]    sboxRom_112;
  wire       [7:0]    sboxRom_113;
  wire       [7:0]    sboxRom_114;
  wire       [7:0]    sboxRom_115;
  wire       [7:0]    sboxRom_116;
  wire       [7:0]    sboxRom_117;
  wire       [7:0]    sboxRom_118;
  wire       [7:0]    sboxRom_119;
  wire       [7:0]    sboxRom_120;
  wire       [7:0]    sboxRom_121;
  wire       [7:0]    sboxRom_122;
  wire       [7:0]    sboxRom_123;
  wire       [7:0]    sboxRom_124;
  wire       [7:0]    sboxRom_125;
  wire       [7:0]    sboxRom_126;
  wire       [7:0]    sboxRom_127;
  wire       [7:0]    sboxRom_128;
  wire       [7:0]    sboxRom_129;
  wire       [7:0]    sboxRom_130;
  wire       [7:0]    sboxRom_131;
  wire       [7:0]    sboxRom_132;
  wire       [7:0]    sboxRom_133;
  wire       [7:0]    sboxRom_134;
  wire       [7:0]    sboxRom_135;
  wire       [7:0]    sboxRom_136;
  wire       [7:0]    sboxRom_137;
  wire       [7:0]    sboxRom_138;
  wire       [7:0]    sboxRom_139;
  wire       [7:0]    sboxRom_140;
  wire       [7:0]    sboxRom_141;
  wire       [7:0]    sboxRom_142;
  wire       [7:0]    sboxRom_143;
  wire       [7:0]    sboxRom_144;
  wire       [7:0]    sboxRom_145;
  wire       [7:0]    sboxRom_146;
  wire       [7:0]    sboxRom_147;
  wire       [7:0]    sboxRom_148;
  wire       [7:0]    sboxRom_149;
  wire       [7:0]    sboxRom_150;
  wire       [7:0]    sboxRom_151;
  wire       [7:0]    sboxRom_152;
  wire       [7:0]    sboxRom_153;
  wire       [7:0]    sboxRom_154;
  wire       [7:0]    sboxRom_155;
  wire       [7:0]    sboxRom_156;
  wire       [7:0]    sboxRom_157;
  wire       [7:0]    sboxRom_158;
  wire       [7:0]    sboxRom_159;
  wire       [7:0]    sboxRom_160;
  wire       [7:0]    sboxRom_161;
  wire       [7:0]    sboxRom_162;
  wire       [7:0]    sboxRom_163;
  wire       [7:0]    sboxRom_164;
  wire       [7:0]    sboxRom_165;
  wire       [7:0]    sboxRom_166;
  wire       [7:0]    sboxRom_167;
  wire       [7:0]    sboxRom_168;
  wire       [7:0]    sboxRom_169;
  wire       [7:0]    sboxRom_170;
  wire       [7:0]    sboxRom_171;
  wire       [7:0]    sboxRom_172;
  wire       [7:0]    sboxRom_173;
  wire       [7:0]    sboxRom_174;
  wire       [7:0]    sboxRom_175;
  wire       [7:0]    sboxRom_176;
  wire       [7:0]    sboxRom_177;
  wire       [7:0]    sboxRom_178;
  wire       [7:0]    sboxRom_179;
  wire       [7:0]    sboxRom_180;
  wire       [7:0]    sboxRom_181;
  wire       [7:0]    sboxRom_182;
  wire       [7:0]    sboxRom_183;
  wire       [7:0]    sboxRom_184;
  wire       [7:0]    sboxRom_185;
  wire       [7:0]    sboxRom_186;
  wire       [7:0]    sboxRom_187;
  wire       [7:0]    sboxRom_188;
  wire       [7:0]    sboxRom_189;
  wire       [7:0]    sboxRom_190;
  wire       [7:0]    sboxRom_191;
  wire       [7:0]    sboxRom_192;
  wire       [7:0]    sboxRom_193;
  wire       [7:0]    sboxRom_194;
  wire       [7:0]    sboxRom_195;
  wire       [7:0]    sboxRom_196;
  wire       [7:0]    sboxRom_197;
  wire       [7:0]    sboxRom_198;
  wire       [7:0]    sboxRom_199;
  wire       [7:0]    sboxRom_200;
  wire       [7:0]    sboxRom_201;
  wire       [7:0]    sboxRom_202;
  wire       [7:0]    sboxRom_203;
  wire       [7:0]    sboxRom_204;
  wire       [7:0]    sboxRom_205;
  wire       [7:0]    sboxRom_206;
  wire       [7:0]    sboxRom_207;
  wire       [7:0]    sboxRom_208;
  wire       [7:0]    sboxRom_209;
  wire       [7:0]    sboxRom_210;
  wire       [7:0]    sboxRom_211;
  wire       [7:0]    sboxRom_212;
  wire       [7:0]    sboxRom_213;
  wire       [7:0]    sboxRom_214;
  wire       [7:0]    sboxRom_215;
  wire       [7:0]    sboxRom_216;
  wire       [7:0]    sboxRom_217;
  wire       [7:0]    sboxRom_218;
  wire       [7:0]    sboxRom_219;
  wire       [7:0]    sboxRom_220;
  wire       [7:0]    sboxRom_221;
  wire       [7:0]    sboxRom_222;
  wire       [7:0]    sboxRom_223;
  wire       [7:0]    sboxRom_224;
  wire       [7:0]    sboxRom_225;
  wire       [7:0]    sboxRom_226;
  wire       [7:0]    sboxRom_227;
  wire       [7:0]    sboxRom_228;
  wire       [7:0]    sboxRom_229;
  wire       [7:0]    sboxRom_230;
  wire       [7:0]    sboxRom_231;
  wire       [7:0]    sboxRom_232;
  wire       [7:0]    sboxRom_233;
  wire       [7:0]    sboxRom_234;
  wire       [7:0]    sboxRom_235;
  wire       [7:0]    sboxRom_236;
  wire       [7:0]    sboxRom_237;
  wire       [7:0]    sboxRom_238;
  wire       [7:0]    sboxRom_239;
  wire       [7:0]    sboxRom_240;
  wire       [7:0]    sboxRom_241;
  wire       [7:0]    sboxRom_242;
  wire       [7:0]    sboxRom_243;
  wire       [7:0]    sboxRom_244;
  wire       [7:0]    sboxRom_245;
  wire       [7:0]    sboxRom_246;
  wire       [7:0]    sboxRom_247;
  wire       [7:0]    sboxRom_248;
  wire       [7:0]    sboxRom_249;
  wire       [7:0]    sboxRom_250;
  wire       [7:0]    sboxRom_251;
  wire       [7:0]    sboxRom_252;
  wire       [7:0]    sboxRom_253;
  wire       [7:0]    sboxRom_254;
  wire       [7:0]    sboxRom_255;
  reg        [127:0]  stateReg;
  reg        [31:0]   roundKeyReg_0;
  reg        [31:0]   roundKeyReg_1;
  reg        [31:0]   roundKeyReg_2;
  reg        [31:0]   roundKeyReg_3;
  reg        [3:0]    roundCount;
  reg                 running;
  reg        [3:0]    rconCounter;
  wire       [7:0]    invSboxRom_0;
  wire       [7:0]    invSboxRom_1;
  wire       [7:0]    invSboxRom_2;
  wire       [7:0]    invSboxRom_3;
  wire       [7:0]    invSboxRom_4;
  wire       [7:0]    invSboxRom_5;
  wire       [7:0]    invSboxRom_6;
  wire       [7:0]    invSboxRom_7;
  wire       [7:0]    invSboxRom_8;
  wire       [7:0]    invSboxRom_9;
  wire       [7:0]    invSboxRom_10;
  wire       [7:0]    invSboxRom_11;
  wire       [7:0]    invSboxRom_12;
  wire       [7:0]    invSboxRom_13;
  wire       [7:0]    invSboxRom_14;
  wire       [7:0]    invSboxRom_15;
  wire       [7:0]    invSboxRom_16;
  wire       [7:0]    invSboxRom_17;
  wire       [7:0]    invSboxRom_18;
  wire       [7:0]    invSboxRom_19;
  wire       [7:0]    invSboxRom_20;
  wire       [7:0]    invSboxRom_21;
  wire       [7:0]    invSboxRom_22;
  wire       [7:0]    invSboxRom_23;
  wire       [7:0]    invSboxRom_24;
  wire       [7:0]    invSboxRom_25;
  wire       [7:0]    invSboxRom_26;
  wire       [7:0]    invSboxRom_27;
  wire       [7:0]    invSboxRom_28;
  wire       [7:0]    invSboxRom_29;
  wire       [7:0]    invSboxRom_30;
  wire       [7:0]    invSboxRom_31;
  wire       [7:0]    invSboxRom_32;
  wire       [7:0]    invSboxRom_33;
  wire       [7:0]    invSboxRom_34;
  wire       [7:0]    invSboxRom_35;
  wire       [7:0]    invSboxRom_36;
  wire       [7:0]    invSboxRom_37;
  wire       [7:0]    invSboxRom_38;
  wire       [7:0]    invSboxRom_39;
  wire       [7:0]    invSboxRom_40;
  wire       [7:0]    invSboxRom_41;
  wire       [7:0]    invSboxRom_42;
  wire       [7:0]    invSboxRom_43;
  wire       [7:0]    invSboxRom_44;
  wire       [7:0]    invSboxRom_45;
  wire       [7:0]    invSboxRom_46;
  wire       [7:0]    invSboxRom_47;
  wire       [7:0]    invSboxRom_48;
  wire       [7:0]    invSboxRom_49;
  wire       [7:0]    invSboxRom_50;
  wire       [7:0]    invSboxRom_51;
  wire       [7:0]    invSboxRom_52;
  wire       [7:0]    invSboxRom_53;
  wire       [7:0]    invSboxRom_54;
  wire       [7:0]    invSboxRom_55;
  wire       [7:0]    invSboxRom_56;
  wire       [7:0]    invSboxRom_57;
  wire       [7:0]    invSboxRom_58;
  wire       [7:0]    invSboxRom_59;
  wire       [7:0]    invSboxRom_60;
  wire       [7:0]    invSboxRom_61;
  wire       [7:0]    invSboxRom_62;
  wire       [7:0]    invSboxRom_63;
  wire       [7:0]    invSboxRom_64;
  wire       [7:0]    invSboxRom_65;
  wire       [7:0]    invSboxRom_66;
  wire       [7:0]    invSboxRom_67;
  wire       [7:0]    invSboxRom_68;
  wire       [7:0]    invSboxRom_69;
  wire       [7:0]    invSboxRom_70;
  wire       [7:0]    invSboxRom_71;
  wire       [7:0]    invSboxRom_72;
  wire       [7:0]    invSboxRom_73;
  wire       [7:0]    invSboxRom_74;
  wire       [7:0]    invSboxRom_75;
  wire       [7:0]    invSboxRom_76;
  wire       [7:0]    invSboxRom_77;
  wire       [7:0]    invSboxRom_78;
  wire       [7:0]    invSboxRom_79;
  wire       [7:0]    invSboxRom_80;
  wire       [7:0]    invSboxRom_81;
  wire       [7:0]    invSboxRom_82;
  wire       [7:0]    invSboxRom_83;
  wire       [7:0]    invSboxRom_84;
  wire       [7:0]    invSboxRom_85;
  wire       [7:0]    invSboxRom_86;
  wire       [7:0]    invSboxRom_87;
  wire       [7:0]    invSboxRom_88;
  wire       [7:0]    invSboxRom_89;
  wire       [7:0]    invSboxRom_90;
  wire       [7:0]    invSboxRom_91;
  wire       [7:0]    invSboxRom_92;
  wire       [7:0]    invSboxRom_93;
  wire       [7:0]    invSboxRom_94;
  wire       [7:0]    invSboxRom_95;
  wire       [7:0]    invSboxRom_96;
  wire       [7:0]    invSboxRom_97;
  wire       [7:0]    invSboxRom_98;
  wire       [7:0]    invSboxRom_99;
  wire       [7:0]    invSboxRom_100;
  wire       [7:0]    invSboxRom_101;
  wire       [7:0]    invSboxRom_102;
  wire       [7:0]    invSboxRom_103;
  wire       [7:0]    invSboxRom_104;
  wire       [7:0]    invSboxRom_105;
  wire       [7:0]    invSboxRom_106;
  wire       [7:0]    invSboxRom_107;
  wire       [7:0]    invSboxRom_108;
  wire       [7:0]    invSboxRom_109;
  wire       [7:0]    invSboxRom_110;
  wire       [7:0]    invSboxRom_111;
  wire       [7:0]    invSboxRom_112;
  wire       [7:0]    invSboxRom_113;
  wire       [7:0]    invSboxRom_114;
  wire       [7:0]    invSboxRom_115;
  wire       [7:0]    invSboxRom_116;
  wire       [7:0]    invSboxRom_117;
  wire       [7:0]    invSboxRom_118;
  wire       [7:0]    invSboxRom_119;
  wire       [7:0]    invSboxRom_120;
  wire       [7:0]    invSboxRom_121;
  wire       [7:0]    invSboxRom_122;
  wire       [7:0]    invSboxRom_123;
  wire       [7:0]    invSboxRom_124;
  wire       [7:0]    invSboxRom_125;
  wire       [7:0]    invSboxRom_126;
  wire       [7:0]    invSboxRom_127;
  wire       [7:0]    invSboxRom_128;
  wire       [7:0]    invSboxRom_129;
  wire       [7:0]    invSboxRom_130;
  wire       [7:0]    invSboxRom_131;
  wire       [7:0]    invSboxRom_132;
  wire       [7:0]    invSboxRom_133;
  wire       [7:0]    invSboxRom_134;
  wire       [7:0]    invSboxRom_135;
  wire       [7:0]    invSboxRom_136;
  wire       [7:0]    invSboxRom_137;
  wire       [7:0]    invSboxRom_138;
  wire       [7:0]    invSboxRom_139;
  wire       [7:0]    invSboxRom_140;
  wire       [7:0]    invSboxRom_141;
  wire       [7:0]    invSboxRom_142;
  wire       [7:0]    invSboxRom_143;
  wire       [7:0]    invSboxRom_144;
  wire       [7:0]    invSboxRom_145;
  wire       [7:0]    invSboxRom_146;
  wire       [7:0]    invSboxRom_147;
  wire       [7:0]    invSboxRom_148;
  wire       [7:0]    invSboxRom_149;
  wire       [7:0]    invSboxRom_150;
  wire       [7:0]    invSboxRom_151;
  wire       [7:0]    invSboxRom_152;
  wire       [7:0]    invSboxRom_153;
  wire       [7:0]    invSboxRom_154;
  wire       [7:0]    invSboxRom_155;
  wire       [7:0]    invSboxRom_156;
  wire       [7:0]    invSboxRom_157;
  wire       [7:0]    invSboxRom_158;
  wire       [7:0]    invSboxRom_159;
  wire       [7:0]    invSboxRom_160;
  wire       [7:0]    invSboxRom_161;
  wire       [7:0]    invSboxRom_162;
  wire       [7:0]    invSboxRom_163;
  wire       [7:0]    invSboxRom_164;
  wire       [7:0]    invSboxRom_165;
  wire       [7:0]    invSboxRom_166;
  wire       [7:0]    invSboxRom_167;
  wire       [7:0]    invSboxRom_168;
  wire       [7:0]    invSboxRom_169;
  wire       [7:0]    invSboxRom_170;
  wire       [7:0]    invSboxRom_171;
  wire       [7:0]    invSboxRom_172;
  wire       [7:0]    invSboxRom_173;
  wire       [7:0]    invSboxRom_174;
  wire       [7:0]    invSboxRom_175;
  wire       [7:0]    invSboxRom_176;
  wire       [7:0]    invSboxRom_177;
  wire       [7:0]    invSboxRom_178;
  wire       [7:0]    invSboxRom_179;
  wire       [7:0]    invSboxRom_180;
  wire       [7:0]    invSboxRom_181;
  wire       [7:0]    invSboxRom_182;
  wire       [7:0]    invSboxRom_183;
  wire       [7:0]    invSboxRom_184;
  wire       [7:0]    invSboxRom_185;
  wire       [7:0]    invSboxRom_186;
  wire       [7:0]    invSboxRom_187;
  wire       [7:0]    invSboxRom_188;
  wire       [7:0]    invSboxRom_189;
  wire       [7:0]    invSboxRom_190;
  wire       [7:0]    invSboxRom_191;
  wire       [7:0]    invSboxRom_192;
  wire       [7:0]    invSboxRom_193;
  wire       [7:0]    invSboxRom_194;
  wire       [7:0]    invSboxRom_195;
  wire       [7:0]    invSboxRom_196;
  wire       [7:0]    invSboxRom_197;
  wire       [7:0]    invSboxRom_198;
  wire       [7:0]    invSboxRom_199;
  wire       [7:0]    invSboxRom_200;
  wire       [7:0]    invSboxRom_201;
  wire       [7:0]    invSboxRom_202;
  wire       [7:0]    invSboxRom_203;
  wire       [7:0]    invSboxRom_204;
  wire       [7:0]    invSboxRom_205;
  wire       [7:0]    invSboxRom_206;
  wire       [7:0]    invSboxRom_207;
  wire       [7:0]    invSboxRom_208;
  wire       [7:0]    invSboxRom_209;
  wire       [7:0]    invSboxRom_210;
  wire       [7:0]    invSboxRom_211;
  wire       [7:0]    invSboxRom_212;
  wire       [7:0]    invSboxRom_213;
  wire       [7:0]    invSboxRom_214;
  wire       [7:0]    invSboxRom_215;
  wire       [7:0]    invSboxRom_216;
  wire       [7:0]    invSboxRom_217;
  wire       [7:0]    invSboxRom_218;
  wire       [7:0]    invSboxRom_219;
  wire       [7:0]    invSboxRom_220;
  wire       [7:0]    invSboxRom_221;
  wire       [7:0]    invSboxRom_222;
  wire       [7:0]    invSboxRom_223;
  wire       [7:0]    invSboxRom_224;
  wire       [7:0]    invSboxRom_225;
  wire       [7:0]    invSboxRom_226;
  wire       [7:0]    invSboxRom_227;
  wire       [7:0]    invSboxRom_228;
  wire       [7:0]    invSboxRom_229;
  wire       [7:0]    invSboxRom_230;
  wire       [7:0]    invSboxRom_231;
  wire       [7:0]    invSboxRom_232;
  wire       [7:0]    invSboxRom_233;
  wire       [7:0]    invSboxRom_234;
  wire       [7:0]    invSboxRom_235;
  wire       [7:0]    invSboxRom_236;
  wire       [7:0]    invSboxRom_237;
  wire       [7:0]    invSboxRom_238;
  wire       [7:0]    invSboxRom_239;
  wire       [7:0]    invSboxRom_240;
  wire       [7:0]    invSboxRom_241;
  wire       [7:0]    invSboxRom_242;
  wire       [7:0]    invSboxRom_243;
  wire       [7:0]    invSboxRom_244;
  wire       [7:0]    invSboxRom_245;
  wire       [7:0]    invSboxRom_246;
  wire       [7:0]    invSboxRom_247;
  wire       [7:0]    invSboxRom_248;
  wire       [7:0]    invSboxRom_249;
  wire       [7:0]    invSboxRom_250;
  wire       [7:0]    invSboxRom_251;
  wire       [7:0]    invSboxRom_252;
  wire       [7:0]    invSboxRom_253;
  wire       [7:0]    invSboxRom_254;
  wire       [7:0]    invSboxRom_255;
  reg                 precomputeRunning;
  reg        [3:0]    precomputeCounter;
  reg        [127:0]  newStateComb;
  reg        [127:0]  rkBitsUsedComb;
  wire                when_AES128_l215;
  wire       [31:0]   _zz_stateReg;
  wire       [31:0]   _zz_stateReg_1;
  wire       [31:0]   _zz_stateReg_2;
  wire       [31:0]   _zz_stateReg_3;
  wire       [7:0]    _zz_stateReg_4;
  wire       [7:0]    _zz_stateReg_5;
  wire       [7:0]    _zz_stateReg_6;
  wire       [7:0]    _zz_stateReg_7;
  wire       [7:0]    _zz_stateReg_8;
  wire       [7:0]    _zz_stateReg_9;
  wire       [7:0]    _zz_stateReg_10;
  wire       [7:0]    _zz_stateReg_11;
  wire       [7:0]    _zz_stateReg_12;
  wire       [7:0]    _zz_stateReg_13;
  wire       [7:0]    _zz_stateReg_14;
  wire       [7:0]    _zz_stateReg_15;
  wire       [7:0]    _zz_stateReg_16;
  wire       [7:0]    _zz_stateReg_17;
  wire       [7:0]    _zz_stateReg_18;
  wire       [7:0]    _zz_stateReg_19;
  reg        [7:0]    _zz_stateReg_20;
  reg        [7:0]    _zz_stateReg_21;
  reg        [7:0]    _zz_stateReg_22;
  reg        [7:0]    _zz_stateReg_23;
  reg        [7:0]    _zz_stateReg_24;
  reg        [7:0]    _zz_stateReg_25;
  reg        [7:0]    _zz_stateReg_26;
  reg        [7:0]    _zz_stateReg_27;
  reg        [7:0]    _zz_stateReg_28;
  reg        [7:0]    _zz_stateReg_29;
  reg        [7:0]    _zz_stateReg_30;
  reg        [7:0]    _zz_stateReg_31;
  reg        [7:0]    _zz_stateReg_32;
  reg        [7:0]    _zz_stateReg_33;
  reg        [7:0]    _zz_stateReg_34;
  reg        [7:0]    _zz_stateReg_35;
  wire                when_AES128_l257;
  wire       [7:0]    _zz_stateReg_36;
  wire       [7:0]    _zz_stateReg_37;
  wire       [7:0]    _zz_stateReg_38;
  wire       [7:0]    _zz_stateReg_39;
  wire       [7:0]    _zz_stateReg_40;
  wire       [7:0]    _zz_stateReg_41;
  wire       [7:0]    _zz_stateReg_42;
  wire       [7:0]    _zz_stateReg_43;
  wire       [7:0]    _zz_stateReg_44;
  wire       [7:0]    _zz_stateReg_45;
  wire       [7:0]    _zz_stateReg_46;
  wire       [7:0]    _zz_stateReg_47;
  wire       [7:0]    _zz_stateReg_48;
  wire       [7:0]    _zz_stateReg_49;
  wire       [7:0]    _zz_stateReg_50;
  wire       [7:0]    _zz_stateReg_51;
  wire       [7:0]    _zz_stateReg_52;
  wire       [7:0]    _zz_stateReg_53;
  wire       [7:0]    _zz_stateReg_54;
  wire       [7:0]    _zz_stateReg_55;
  wire       [7:0]    _zz_stateReg_56;
  wire       [7:0]    _zz_stateReg_57;
  wire       [7:0]    _zz_stateReg_58;
  wire       [7:0]    _zz_stateReg_59;
  wire       [7:0]    _zz_stateReg_60;
  wire       [7:0]    _zz_stateReg_61;
  wire       [7:0]    _zz_stateReg_62;
  wire       [7:0]    _zz_stateReg_63;
  wire       [7:0]    _zz_stateReg_64;
  wire       [7:0]    _zz_stateReg_65;
  wire       [7:0]    _zz_stateReg_66;
  wire       [7:0]    _zz_stateReg_67;
  wire       [127:0]  _zz_stateReg_68;
  wire       [7:0]    _zz_roundKeyReg_0;
  wire       [31:0]   _zz_roundKeyReg_0_1;
  wire       [31:0]   _zz_roundKeyReg_0_2;
  wire       [31:0]   _zz_roundKeyReg_1;
  wire       [31:0]   _zz_roundKeyReg_2;
  wire       [31:0]   _zz_roundKeyReg_3;
  wire       [127:0]  _zz_stateReg_69;
  wire                when_AES128_l291;
  wire                when_AES128_l297;
  wire       [31:0]   _zz_stateReg_70;
  wire       [31:0]   _zz_stateReg_71;
  wire       [31:0]   _zz_stateReg_72;
  wire       [31:0]   _zz_stateReg_73;
  wire       [31:0]   _zz_stateReg_74;
  wire                when_AES128_l313;
  wire       [31:0]   _zz_roundKeyReg_3_1;
  wire       [31:0]   _zz_roundKeyReg_2_1;
  wire       [31:0]   _zz_roundKeyReg_1_1;
  wire       [31:0]   _zz_roundKeyReg_0_3;
  wire       [31:0]   _zz_roundKeyReg_0_4;
  wire       [127:0]  _zz_stateReg_75;
  wire       [7:0]    _zz_stateReg_76;
  wire       [7:0]    _zz_stateReg_77;
  wire       [7:0]    _zz_stateReg_78;
  wire       [7:0]    _zz_stateReg_79;
  wire       [7:0]    _zz_stateReg_80;
  wire       [7:0]    _zz_stateReg_81;
  wire       [7:0]    _zz_stateReg_82;
  wire       [7:0]    _zz_stateReg_83;
  wire       [7:0]    _zz_stateReg_84;
  wire       [7:0]    _zz_stateReg_85;
  wire       [7:0]    _zz_stateReg_86;
  wire       [7:0]    _zz_stateReg_87;
  wire       [7:0]    _zz_stateReg_88;
  wire       [7:0]    _zz_stateReg_89;
  wire       [7:0]    _zz_stateReg_90;
  wire       [7:0]    _zz_stateReg_91;
  reg        [7:0]    _zz_stateReg_92;
  reg        [7:0]    _zz_stateReg_93;
  reg        [7:0]    _zz_stateReg_94;
  reg        [7:0]    _zz_stateReg_95;
  reg        [7:0]    _zz_stateReg_96;
  reg        [7:0]    _zz_stateReg_97;
  reg        [7:0]    _zz_stateReg_98;
  reg        [7:0]    _zz_stateReg_99;
  reg        [7:0]    _zz_stateReg_100;
  reg        [7:0]    _zz_stateReg_101;
  reg        [7:0]    _zz_stateReg_102;
  reg        [7:0]    _zz_stateReg_103;
  reg        [7:0]    _zz_stateReg_104;
  reg        [7:0]    _zz_stateReg_105;
  reg        [7:0]    _zz_stateReg_106;
  reg        [7:0]    _zz_stateReg_107;
  wire                when_AES128_l356;
  wire       [7:0]    _zz_stateReg_108;
  wire       [7:0]    _zz_stateReg_109;
  wire       [7:0]    _zz_stateReg_110;
  wire       [7:0]    _zz_stateReg_111;
  wire       [7:0]    _zz_stateReg_112;
  wire       [7:0]    _zz_stateReg_113;
  wire       [7:0]    _zz_stateReg_114;
  wire       [7:0]    _zz_stateReg_115;
  wire       [7:0]    _zz_stateReg_116;
  wire       [7:0]    _zz_stateReg_117;
  wire       [7:0]    _zz_stateReg_118;
  wire       [7:0]    _zz_stateReg_119;
  wire       [7:0]    _zz_stateReg_120;
  wire       [7:0]    _zz_stateReg_121;
  wire       [7:0]    _zz_stateReg_122;
  wire       [7:0]    _zz_stateReg_123;
  wire       [7:0]    _zz_stateReg_124;
  wire       [7:0]    _zz_stateReg_125;
  wire       [7:0]    _zz_stateReg_126;
  wire       [7:0]    _zz_stateReg_127;
  wire       [7:0]    _zz_stateReg_128;
  wire       [7:0]    _zz_stateReg_129;
  wire       [7:0]    _zz_stateReg_130;
  wire       [7:0]    _zz_stateReg_131;
  wire       [7:0]    _zz_stateReg_132;
  wire       [7:0]    _zz_stateReg_133;
  wire       [7:0]    _zz_stateReg_134;
  wire       [7:0]    _zz_stateReg_135;
  wire       [7:0]    _zz_stateReg_136;
  wire       [7:0]    _zz_stateReg_137;
  wire       [7:0]    _zz_stateReg_138;
  wire       [7:0]    _zz_stateReg_139;
  wire       [7:0]    _zz_stateReg_140;
  wire       [7:0]    _zz_stateReg_141;
  wire       [7:0]    _zz_stateReg_142;
  wire       [7:0]    _zz_stateReg_143;
  wire       [7:0]    _zz_stateReg_144;
  wire       [7:0]    _zz_stateReg_145;
  wire       [7:0]    _zz_stateReg_146;
  wire       [7:0]    _zz_stateReg_147;
  wire       [7:0]    _zz_stateReg_148;
  wire       [7:0]    _zz_stateReg_149;
  wire       [7:0]    _zz_stateReg_150;
  wire       [7:0]    _zz_stateReg_151;
  wire       [7:0]    _zz_stateReg_152;
  wire       [7:0]    _zz_stateReg_153;
  wire       [7:0]    _zz_stateReg_154;
  wire       [7:0]    _zz_stateReg_155;
  wire       [7:0]    _zz_stateReg_156;
  wire       [7:0]    _zz_stateReg_157;
  wire       [7:0]    _zz_stateReg_158;
  wire       [7:0]    _zz_stateReg_159;
  wire       [7:0]    _zz_stateReg_160;
  wire       [7:0]    _zz_stateReg_161;
  wire       [7:0]    _zz_stateReg_162;
  wire       [7:0]    _zz_stateReg_163;
  wire       [7:0]    _zz_stateReg_164;
  wire       [7:0]    _zz_stateReg_165;
  wire       [7:0]    _zz_stateReg_166;
  wire       [7:0]    _zz_stateReg_167;
  wire       [7:0]    _zz_stateReg_168;
  wire       [7:0]    _zz_stateReg_169;
  wire       [7:0]    _zz_stateReg_170;
  wire       [7:0]    _zz_stateReg_171;
  wire       [7:0]    _zz_stateReg_172;
  wire       [7:0]    _zz_stateReg_173;
  wire       [7:0]    _zz_stateReg_174;
  wire       [7:0]    _zz_stateReg_175;
  wire       [7:0]    _zz_stateReg_176;
  wire       [7:0]    _zz_stateReg_177;
  wire       [7:0]    _zz_stateReg_178;
  wire       [7:0]    _zz_stateReg_179;
  wire       [7:0]    _zz_stateReg_180;
  wire       [7:0]    _zz_stateReg_181;
  wire       [7:0]    _zz_stateReg_182;
  wire       [7:0]    _zz_stateReg_183;
  wire       [7:0]    _zz_stateReg_184;
  wire       [7:0]    _zz_stateReg_185;
  wire       [7:0]    _zz_stateReg_186;
  wire       [7:0]    _zz_stateReg_187;
  wire       [7:0]    _zz_stateReg_188;
  wire       [7:0]    _zz_stateReg_189;
  wire       [7:0]    _zz_stateReg_190;
  wire       [7:0]    _zz_stateReg_191;
  wire       [7:0]    _zz_stateReg_192;
  wire       [7:0]    _zz_stateReg_193;
  wire       [7:0]    _zz_stateReg_194;
  wire       [7:0]    _zz_stateReg_195;
  wire       [7:0]    _zz_stateReg_196;
  wire       [7:0]    _zz_stateReg_197;
  wire       [7:0]    _zz_stateReg_198;
  wire       [7:0]    _zz_stateReg_199;
  wire       [7:0]    _zz_stateReg_200;
  wire       [7:0]    _zz_stateReg_201;
  wire       [7:0]    _zz_stateReg_202;
  wire       [7:0]    _zz_stateReg_203;
  wire       [7:0]    _zz_stateReg_204;
  wire       [7:0]    _zz_stateReg_205;
  wire       [7:0]    _zz_stateReg_206;
  wire       [7:0]    _zz_stateReg_207;
  wire       [7:0]    _zz_stateReg_208;
  wire       [7:0]    _zz_stateReg_209;
  wire       [7:0]    _zz_stateReg_210;
  wire       [7:0]    _zz_stateReg_211;
  wire       [7:0]    _zz_stateReg_212;
  wire       [7:0]    _zz_stateReg_213;
  wire       [7:0]    _zz_stateReg_214;
  wire       [7:0]    _zz_stateReg_215;
  wire       [7:0]    _zz_stateReg_216;
  wire       [7:0]    _zz_stateReg_217;
  wire       [7:0]    _zz_stateReg_218;
  wire       [7:0]    _zz_stateReg_219;
  wire       [7:0]    _zz_stateReg_220;
  wire       [7:0]    _zz_stateReg_221;
  wire       [7:0]    _zz_stateReg_222;
  wire       [7:0]    _zz_stateReg_223;
  wire       [7:0]    _zz_stateReg_224;
  wire       [7:0]    _zz_stateReg_225;
  wire       [7:0]    _zz_stateReg_226;
  wire       [7:0]    _zz_stateReg_227;
  wire       [7:0]    _zz_stateReg_228;
  wire       [7:0]    _zz_stateReg_229;
  wire       [7:0]    _zz_stateReg_230;
  wire       [7:0]    _zz_stateReg_231;
  wire       [7:0]    _zz_stateReg_232;
  wire       [7:0]    _zz_stateReg_233;
  wire       [7:0]    _zz_stateReg_234;
  wire       [7:0]    _zz_stateReg_235;
  wire       [7:0]    _zz_stateReg_236;
  wire       [7:0]    _zz_stateReg_237;
  wire       [7:0]    _zz_stateReg_238;
  wire       [7:0]    _zz_stateReg_239;
  wire       [7:0]    _zz_stateReg_240;
  wire       [7:0]    _zz_stateReg_241;
  wire       [7:0]    _zz_stateReg_242;
  wire       [7:0]    _zz_stateReg_243;
  wire       [7:0]    _zz_stateReg_244;
  wire       [7:0]    _zz_stateReg_245;
  wire       [7:0]    _zz_stateReg_246;
  wire       [7:0]    _zz_stateReg_247;
  wire       [7:0]    _zz_stateReg_248;
  wire       [7:0]    _zz_stateReg_249;
  wire       [7:0]    _zz_stateReg_250;
  wire       [7:0]    _zz_stateReg_251;
  wire       [7:0]    _zz_stateReg_252;
  wire       [7:0]    _zz_stateReg_253;
  wire       [7:0]    _zz_stateReg_254;
  wire       [7:0]    _zz_stateReg_255;
  wire       [7:0]    _zz_stateReg_256;
  wire       [7:0]    _zz_stateReg_257;
  wire       [7:0]    _zz_stateReg_258;
  wire       [7:0]    _zz_stateReg_259;
  wire       [7:0]    _zz_stateReg_260;
  wire       [7:0]    _zz_stateReg_261;
  wire       [7:0]    _zz_stateReg_262;
  wire       [7:0]    _zz_stateReg_263;
  wire       [7:0]    _zz_stateReg_264;
  wire       [7:0]    _zz_stateReg_265;
  wire       [7:0]    _zz_stateReg_266;
  wire       [7:0]    _zz_stateReg_267;
  wire       [7:0]    _zz_stateReg_268;
  wire       [7:0]    _zz_stateReg_269;
  wire       [7:0]    _zz_stateReg_270;
  wire       [7:0]    _zz_stateReg_271;
  wire       [7:0]    _zz_stateReg_272;
  wire       [7:0]    _zz_stateReg_273;
  wire       [7:0]    _zz_stateReg_274;
  wire       [7:0]    _zz_stateReg_275;
  wire       [7:0]    _zz_stateReg_276;
  wire       [7:0]    _zz_stateReg_277;
  wire       [7:0]    _zz_stateReg_278;
  wire       [7:0]    _zz_stateReg_279;
  wire       [7:0]    _zz_stateReg_280;
  wire       [7:0]    _zz_stateReg_281;
  wire       [7:0]    _zz_stateReg_282;
  wire       [7:0]    _zz_stateReg_283;
  wire       [7:0]    _zz_stateReg_284;
  wire       [7:0]    _zz_stateReg_285;
  wire       [7:0]    _zz_stateReg_286;
  wire       [7:0]    _zz_stateReg_287;
  wire       [7:0]    _zz_stateReg_288;
  wire       [7:0]    _zz_stateReg_289;
  wire       [7:0]    _zz_stateReg_290;
  wire       [7:0]    _zz_stateReg_291;
  wire       [7:0]    _zz_stateReg_292;
  wire       [7:0]    _zz_stateReg_293;
  wire       [7:0]    _zz_stateReg_294;
  wire       [7:0]    _zz_stateReg_295;
  wire       [7:0]    _zz_stateReg_296;
  wire       [7:0]    _zz_stateReg_297;
  wire       [7:0]    _zz_stateReg_298;
  wire       [7:0]    _zz_stateReg_299;
  wire       [7:0]    _zz_stateReg_300;
  wire       [7:0]    _zz_stateReg_301;
  wire       [7:0]    _zz_stateReg_302;
  wire       [7:0]    _zz_stateReg_303;
  wire       [7:0]    _zz_stateReg_304;
  wire       [7:0]    _zz_stateReg_305;
  wire       [7:0]    _zz_stateReg_306;
  wire       [7:0]    _zz_stateReg_307;
  wire       [7:0]    _zz_stateReg_308;
  wire       [7:0]    _zz_stateReg_309;
  wire       [7:0]    _zz_stateReg_310;
  wire       [7:0]    _zz_stateReg_311;
  wire       [7:0]    _zz_stateReg_312;
  wire       [7:0]    _zz_stateReg_313;
  wire       [7:0]    _zz_stateReg_314;
  wire       [7:0]    _zz_stateReg_315;
  wire       [7:0]    _zz_stateReg_316;
  wire       [7:0]    _zz_stateReg_317;
  wire       [7:0]    _zz_stateReg_318;
  wire       [7:0]    _zz_stateReg_319;
  wire       [7:0]    _zz_stateReg_320;
  wire       [7:0]    _zz_stateReg_321;
  wire       [7:0]    _zz_stateReg_322;
  wire       [7:0]    _zz_stateReg_323;
  wire       [7:0]    _zz_stateReg_324;
  wire       [7:0]    _zz_stateReg_325;
  wire       [7:0]    _zz_stateReg_326;
  wire       [7:0]    _zz_stateReg_327;
  wire       [7:0]    _zz_stateReg_328;
  wire       [7:0]    _zz_stateReg_329;
  wire       [7:0]    _zz_stateReg_330;
  wire       [7:0]    _zz_stateReg_331;
  wire       [7:0]    _zz_stateReg_332;
  wire       [7:0]    _zz_stateReg_333;
  wire       [7:0]    _zz_stateReg_334;
  wire       [7:0]    _zz_stateReg_335;
  wire       [7:0]    _zz_stateReg_336;
  wire       [7:0]    _zz_stateReg_337;
  wire       [7:0]    _zz_stateReg_338;
  wire       [7:0]    _zz_stateReg_339;
  wire       [7:0]    _zz_stateReg_340;
  wire       [7:0]    _zz_stateReg_341;
  wire       [7:0]    _zz_stateReg_342;
  wire       [7:0]    _zz_stateReg_343;
  wire       [7:0]    _zz_stateReg_344;
  wire       [7:0]    _zz_stateReg_345;
  wire       [7:0]    _zz_stateReg_346;
  wire       [7:0]    _zz_stateReg_347;
  wire       [7:0]    _zz_stateReg_348;
  wire       [7:0]    _zz_stateReg_349;
  wire       [7:0]    _zz_stateReg_350;
  wire       [7:0]    _zz_stateReg_351;
  wire       [7:0]    _zz_stateReg_352;
  wire       [7:0]    _zz_stateReg_353;
  wire       [7:0]    _zz_stateReg_354;
  wire       [7:0]    _zz_stateReg_355;
  wire       [7:0]    _zz_stateReg_356;
  wire       [7:0]    _zz_stateReg_357;
  wire       [7:0]    _zz_stateReg_358;
  wire       [7:0]    _zz_stateReg_359;
  wire       [7:0]    _zz_stateReg_360;
  wire       [7:0]    _zz_stateReg_361;
  wire       [7:0]    _zz_stateReg_362;
  wire       [7:0]    _zz_stateReg_363;
  wire       [7:0]    _zz_stateReg_364;
  wire       [7:0]    _zz_stateReg_365;
  wire       [7:0]    _zz_stateReg_366;
  wire       [7:0]    _zz_stateReg_367;
  wire       [7:0]    _zz_stateReg_368;
  wire       [7:0]    _zz_stateReg_369;
  wire       [7:0]    _zz_stateReg_370;
  wire       [7:0]    _zz_stateReg_371;
  wire       [7:0]    _zz_stateReg_372;
  wire       [7:0]    _zz_stateReg_373;
  wire       [7:0]    _zz_stateReg_374;
  wire       [7:0]    _zz_stateReg_375;
  wire       [7:0]    _zz_stateReg_376;
  wire       [7:0]    _zz_stateReg_377;
  wire       [7:0]    _zz_stateReg_378;
  wire       [7:0]    _zz_stateReg_379;
  wire       [7:0]    _zz_stateReg_380;
  wire       [7:0]    _zz_stateReg_381;
  wire       [7:0]    _zz_stateReg_382;
  wire       [7:0]    _zz_stateReg_383;
  wire       [7:0]    _zz_stateReg_384;
  wire       [7:0]    _zz_stateReg_385;
  wire       [7:0]    _zz_stateReg_386;
  wire       [7:0]    _zz_stateReg_387;
  wire       [7:0]    _zz_stateReg_388;
  wire       [7:0]    _zz_stateReg_389;
  wire       [7:0]    _zz_stateReg_390;
  wire       [7:0]    _zz_stateReg_391;
  wire       [7:0]    _zz_stateReg_392;
  wire       [7:0]    _zz_stateReg_393;
  wire       [7:0]    _zz_stateReg_394;
  wire       [7:0]    _zz_stateReg_395;
  wire       [7:0]    _zz_stateReg_396;
  wire       [7:0]    _zz_stateReg_397;
  wire       [7:0]    _zz_stateReg_398;
  wire       [7:0]    _zz_stateReg_399;
  wire       [7:0]    _zz_stateReg_400;
  wire       [7:0]    _zz_stateReg_401;
  wire       [7:0]    _zz_stateReg_402;
  wire       [7:0]    _zz_stateReg_403;
  wire       [7:0]    _zz_stateReg_404;
  wire       [7:0]    _zz_stateReg_405;
  wire       [7:0]    _zz_stateReg_406;
  wire       [7:0]    _zz_stateReg_407;
  wire       [7:0]    _zz_stateReg_408;
  wire       [7:0]    _zz_stateReg_409;
  wire       [7:0]    _zz_stateReg_410;
  wire       [7:0]    _zz_stateReg_411;
  wire       [7:0]    _zz_stateReg_412;
  wire       [7:0]    _zz_stateReg_413;
  wire       [7:0]    _zz_stateReg_414;
  wire       [7:0]    _zz_stateReg_415;
  wire       [7:0]    _zz_stateReg_416;
  wire       [7:0]    _zz_stateReg_417;
  wire       [7:0]    _zz_stateReg_418;
  wire       [7:0]    _zz_stateReg_419;
  wire       [7:0]    _zz_stateReg_420;
  wire       [7:0]    _zz_stateReg_421;
  wire       [7:0]    _zz_stateReg_422;
  wire       [7:0]    _zz_stateReg_423;
  wire       [7:0]    _zz_stateReg_424;
  wire       [7:0]    _zz_stateReg_425;
  wire       [7:0]    _zz_stateReg_426;
  wire       [7:0]    _zz_stateReg_427;
  wire       [7:0]    _zz_stateReg_428;
  wire       [7:0]    _zz_stateReg_429;
  wire       [7:0]    _zz_stateReg_430;
  wire       [7:0]    _zz_stateReg_431;
  wire       [7:0]    _zz_stateReg_432;
  wire       [7:0]    _zz_stateReg_433;
  wire       [7:0]    _zz_stateReg_434;
  wire       [7:0]    _zz_stateReg_435;
  wire       [7:0]    _zz_stateReg_436;
  wire       [7:0]    _zz_stateReg_437;
  wire       [7:0]    _zz_stateReg_438;
  wire       [7:0]    _zz_stateReg_439;
  wire       [7:0]    _zz_stateReg_440;
  wire       [7:0]    _zz_stateReg_441;
  wire       [7:0]    _zz_stateReg_442;
  wire       [7:0]    _zz_stateReg_443;
  wire       [7:0]    _zz_stateReg_444;
  wire       [7:0]    _zz_stateReg_445;
  wire       [7:0]    _zz_stateReg_446;
  wire       [7:0]    _zz_stateReg_447;
  wire       [7:0]    _zz_stateReg_448;
  wire       [7:0]    _zz_stateReg_449;
  wire       [7:0]    _zz_stateReg_450;
  wire       [7:0]    _zz_stateReg_451;
  wire       [7:0]    _zz_stateReg_452;
  wire       [7:0]    _zz_stateReg_453;
  wire       [7:0]    _zz_stateReg_454;
  wire       [7:0]    _zz_stateReg_455;
  wire       [7:0]    _zz_stateReg_456;
  wire       [7:0]    _zz_stateReg_457;
  wire       [7:0]    _zz_stateReg_458;
  wire       [7:0]    _zz_stateReg_459;
  wire       [7:0]    _zz_stateReg_460;
  wire       [7:0]    _zz_stateReg_461;
  wire       [7:0]    _zz_stateReg_462;
  wire       [7:0]    _zz_stateReg_463;
  wire       [7:0]    _zz_stateReg_464;
  wire       [7:0]    _zz_stateReg_465;
  wire       [7:0]    _zz_stateReg_466;
  wire       [7:0]    _zz_stateReg_467;
  wire       [7:0]    _zz_stateReg_468;
  wire       [7:0]    _zz_stateReg_469;
  wire       [7:0]    _zz_stateReg_470;
  wire       [7:0]    _zz_stateReg_471;
  wire       [7:0]    _zz_stateReg_472;
  wire       [7:0]    _zz_stateReg_473;
  wire       [7:0]    _zz_stateReg_474;
  wire       [7:0]    _zz_stateReg_475;
  wire       [7:0]    _zz_stateReg_476;
  wire       [7:0]    _zz_stateReg_477;
  wire       [7:0]    _zz_stateReg_478;
  wire       [7:0]    _zz_stateReg_479;
  wire       [7:0]    _zz_stateReg_480;
  wire       [7:0]    _zz_stateReg_481;
  wire       [7:0]    _zz_stateReg_482;
  wire       [7:0]    _zz_stateReg_483;
  wire       [7:0]    _zz_stateReg_484;
  wire       [7:0]    _zz_stateReg_485;
  wire       [7:0]    _zz_stateReg_486;
  wire       [7:0]    _zz_stateReg_487;
  wire       [7:0]    _zz_stateReg_488;
  wire       [7:0]    _zz_stateReg_489;
  wire       [7:0]    _zz_stateReg_490;
  wire       [7:0]    _zz_stateReg_491;
  wire       [7:0]    _zz_stateReg_492;
  wire       [7:0]    _zz_stateReg_493;
  wire       [7:0]    _zz_stateReg_494;
  wire       [7:0]    _zz_stateReg_495;
  wire       [7:0]    _zz_stateReg_496;
  wire       [7:0]    _zz_stateReg_497;
  wire       [7:0]    _zz_stateReg_498;
  wire       [7:0]    _zz_stateReg_499;
  wire       [7:0]    _zz_stateReg_500;
  wire       [7:0]    _zz_stateReg_501;
  wire       [7:0]    _zz_stateReg_502;
  wire       [7:0]    _zz_stateReg_503;
  wire       [7:0]    _zz_stateReg_504;
  wire       [7:0]    _zz_stateReg_505;
  wire       [7:0]    _zz_stateReg_506;
  wire       [7:0]    _zz_stateReg_507;
  wire       [7:0]    _zz_stateReg_508;
  wire       [7:0]    _zz_stateReg_509;
  wire       [7:0]    _zz_stateReg_510;
  wire       [7:0]    _zz_stateReg_511;
  wire       [7:0]    _zz_stateReg_512;
  wire       [7:0]    _zz_stateReg_513;
  wire       [7:0]    _zz_stateReg_514;
  wire       [7:0]    _zz_stateReg_515;
  wire       [7:0]    _zz_stateReg_516;
  wire       [7:0]    _zz_stateReg_517;
  wire       [7:0]    _zz_stateReg_518;
  wire       [7:0]    _zz_stateReg_519;
  wire       [7:0]    _zz_stateReg_520;
  wire       [7:0]    _zz_stateReg_521;
  wire       [7:0]    _zz_stateReg_522;
  wire       [7:0]    _zz_stateReg_523;
  wire       [7:0]    _zz_stateReg_524;
  wire       [7:0]    _zz_stateReg_525;
  wire       [7:0]    _zz_stateReg_526;
  wire       [7:0]    _zz_stateReg_527;
  wire       [7:0]    _zz_stateReg_528;
  wire       [7:0]    _zz_stateReg_529;
  wire       [7:0]    _zz_stateReg_530;
  wire       [7:0]    _zz_stateReg_531;
  wire       [7:0]    _zz_stateReg_532;
  wire       [7:0]    _zz_stateReg_533;
  wire       [7:0]    _zz_stateReg_534;
  wire       [7:0]    _zz_stateReg_535;
  wire       [7:0]    _zz_stateReg_536;
  wire       [7:0]    _zz_stateReg_537;
  wire       [7:0]    _zz_stateReg_538;
  wire       [7:0]    _zz_stateReg_539;
  wire       [7:0]    _zz_stateReg_540;
  wire       [7:0]    _zz_stateReg_541;
  wire       [7:0]    _zz_stateReg_542;
  wire       [7:0]    _zz_stateReg_543;
  wire       [7:0]    _zz_stateReg_544;
  wire       [7:0]    _zz_stateReg_545;
  wire       [7:0]    _zz_stateReg_546;
  wire       [7:0]    _zz_stateReg_547;
  wire       [7:0]    _zz_stateReg_548;
  wire       [7:0]    _zz_stateReg_549;
  wire       [7:0]    _zz_stateReg_550;
  wire       [7:0]    _zz_stateReg_551;
  wire       [7:0]    _zz_stateReg_552;
  wire       [7:0]    _zz_stateReg_553;
  wire       [7:0]    _zz_stateReg_554;
  wire       [7:0]    _zz_stateReg_555;
  wire                when_AES128_l383;
  wire                when_AES128_l389;
  wire                when_AES128_l229;
  wire                when_AES128_l299;
  wire                when_AES128_l324;

  assign _zz__zz_stateReg_36 = ({1'd0,_zz_stateReg_4} <<< 1'd1);
  assign _zz__zz_stateReg_37 = ({1'd0,_zz_stateReg_5} <<< 1'd1);
  assign _zz__zz_stateReg_38 = ({1'd0,_zz_stateReg_5} <<< 1'd1);
  assign _zz__zz_stateReg_39 = ({1'd0,_zz_stateReg_6} <<< 1'd1);
  assign _zz__zz_stateReg_40 = ({1'd0,_zz_stateReg_6} <<< 1'd1);
  assign _zz__zz_stateReg_41 = ({1'd0,_zz_stateReg_7} <<< 1'd1);
  assign _zz__zz_stateReg_42 = ({1'd0,_zz_stateReg_4} <<< 1'd1);
  assign _zz__zz_stateReg_43 = ({1'd0,_zz_stateReg_7} <<< 1'd1);
  assign _zz__zz_stateReg_44 = ({1'd0,_zz_stateReg_8} <<< 1'd1);
  assign _zz__zz_stateReg_45 = ({1'd0,_zz_stateReg_9} <<< 1'd1);
  assign _zz__zz_stateReg_46 = ({1'd0,_zz_stateReg_9} <<< 1'd1);
  assign _zz__zz_stateReg_47 = ({1'd0,_zz_stateReg_10} <<< 1'd1);
  assign _zz__zz_stateReg_48 = ({1'd0,_zz_stateReg_10} <<< 1'd1);
  assign _zz__zz_stateReg_49 = ({1'd0,_zz_stateReg_11} <<< 1'd1);
  assign _zz__zz_stateReg_50 = ({1'd0,_zz_stateReg_8} <<< 1'd1);
  assign _zz__zz_stateReg_51 = ({1'd0,_zz_stateReg_11} <<< 1'd1);
  assign _zz__zz_stateReg_52 = ({1'd0,_zz_stateReg_12} <<< 1'd1);
  assign _zz__zz_stateReg_53 = ({1'd0,_zz_stateReg_13} <<< 1'd1);
  assign _zz__zz_stateReg_54 = ({1'd0,_zz_stateReg_13} <<< 1'd1);
  assign _zz__zz_stateReg_55 = ({1'd0,_zz_stateReg_14} <<< 1'd1);
  assign _zz__zz_stateReg_56 = ({1'd0,_zz_stateReg_14} <<< 1'd1);
  assign _zz__zz_stateReg_57 = ({1'd0,_zz_stateReg_15} <<< 1'd1);
  assign _zz__zz_stateReg_58 = ({1'd0,_zz_stateReg_12} <<< 1'd1);
  assign _zz__zz_stateReg_59 = ({1'd0,_zz_stateReg_15} <<< 1'd1);
  assign _zz__zz_stateReg_60 = ({1'd0,_zz_stateReg_16} <<< 1'd1);
  assign _zz__zz_stateReg_61 = ({1'd0,_zz_stateReg_17} <<< 1'd1);
  assign _zz__zz_stateReg_62 = ({1'd0,_zz_stateReg_17} <<< 1'd1);
  assign _zz__zz_stateReg_63 = ({1'd0,_zz_stateReg_18} <<< 1'd1);
  assign _zz__zz_stateReg_64 = ({1'd0,_zz_stateReg_18} <<< 1'd1);
  assign _zz__zz_stateReg_65 = ({1'd0,_zz_stateReg_19} <<< 1'd1);
  assign _zz__zz_stateReg_66 = ({1'd0,_zz_stateReg_16} <<< 1'd1);
  assign _zz__zz_stateReg_67 = ({1'd0,_zz_stateReg_19} <<< 1'd1);
  assign _zz__zz_stateReg_108 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_110 = ({1'd0,_zz_stateReg_109} <<< 1'd1);
  assign _zz__zz_stateReg_112 = ({1'd0,_zz_stateReg_111} <<< 1'd1);
  assign _zz__zz_stateReg_113 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_115 = ({1'd0,_zz_stateReg_114} <<< 1'd1);
  assign _zz__zz_stateReg_116 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_117 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_119 = ({1'd0,_zz_stateReg_118} <<< 1'd1);
  assign _zz__zz_stateReg_121 = ({1'd0,_zz_stateReg_120} <<< 1'd1);
  assign _zz__zz_stateReg_122 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_123 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_125 = ({1'd0,_zz_stateReg_124} <<< 1'd1);
  assign _zz__zz_stateReg_127 = ({1'd0,_zz_stateReg_126} <<< 1'd1);
  assign _zz__zz_stateReg_128 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_130 = ({1'd0,_zz_stateReg_129} <<< 1'd1);
  assign _zz__zz_stateReg_131 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_133 = ({1'd0,_zz_stateReg_132} <<< 1'd1);
  assign _zz__zz_stateReg_135 = ({1'd0,_zz_stateReg_134} <<< 1'd1);
  assign _zz__zz_stateReg_136 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_138 = ({1'd0,_zz_stateReg_137} <<< 1'd1);
  assign _zz__zz_stateReg_140 = ({1'd0,_zz_stateReg_139} <<< 1'd1);
  assign _zz__zz_stateReg_141 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_143 = ({1'd0,_zz_stateReg_142} <<< 1'd1);
  assign _zz__zz_stateReg_145 = ({1'd0,_zz_stateReg_144} <<< 1'd1);
  assign _zz__zz_stateReg_146 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_148 = ({1'd0,_zz_stateReg_147} <<< 1'd1);
  assign _zz__zz_stateReg_149 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_150 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_152 = ({1'd0,_zz_stateReg_151} <<< 1'd1);
  assign _zz__zz_stateReg_154 = ({1'd0,_zz_stateReg_153} <<< 1'd1);
  assign _zz__zz_stateReg_155 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_156 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_158 = ({1'd0,_zz_stateReg_157} <<< 1'd1);
  assign _zz__zz_stateReg_160 = ({1'd0,_zz_stateReg_159} <<< 1'd1);
  assign _zz__zz_stateReg_161 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_163 = ({1'd0,_zz_stateReg_162} <<< 1'd1);
  assign _zz__zz_stateReg_164 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_166 = ({1'd0,_zz_stateReg_165} <<< 1'd1);
  assign _zz__zz_stateReg_168 = ({1'd0,_zz_stateReg_167} <<< 1'd1);
  assign _zz__zz_stateReg_169 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_171 = ({1'd0,_zz_stateReg_170} <<< 1'd1);
  assign _zz__zz_stateReg_172 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_174 = ({1'd0,_zz_stateReg_173} <<< 1'd1);
  assign _zz__zz_stateReg_176 = ({1'd0,_zz_stateReg_175} <<< 1'd1);
  assign _zz__zz_stateReg_177 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_179 = ({1'd0,_zz_stateReg_178} <<< 1'd1);
  assign _zz__zz_stateReg_181 = ({1'd0,_zz_stateReg_180} <<< 1'd1);
  assign _zz__zz_stateReg_182 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_184 = ({1'd0,_zz_stateReg_183} <<< 1'd1);
  assign _zz__zz_stateReg_185 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_186 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_188 = ({1'd0,_zz_stateReg_187} <<< 1'd1);
  assign _zz__zz_stateReg_190 = ({1'd0,_zz_stateReg_189} <<< 1'd1);
  assign _zz__zz_stateReg_191 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_192 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_194 = ({1'd0,_zz_stateReg_193} <<< 1'd1);
  assign _zz__zz_stateReg_196 = ({1'd0,_zz_stateReg_195} <<< 1'd1);
  assign _zz__zz_stateReg_197 = ({1'd0,_zz_stateReg_76} <<< 1'd1);
  assign _zz__zz_stateReg_198 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_200 = ({1'd0,_zz_stateReg_199} <<< 1'd1);
  assign _zz__zz_stateReg_202 = ({1'd0,_zz_stateReg_201} <<< 1'd1);
  assign _zz__zz_stateReg_203 = ({1'd0,_zz_stateReg_77} <<< 1'd1);
  assign _zz__zz_stateReg_205 = ({1'd0,_zz_stateReg_204} <<< 1'd1);
  assign _zz__zz_stateReg_206 = ({1'd0,_zz_stateReg_78} <<< 1'd1);
  assign _zz__zz_stateReg_208 = ({1'd0,_zz_stateReg_207} <<< 1'd1);
  assign _zz__zz_stateReg_210 = ({1'd0,_zz_stateReg_209} <<< 1'd1);
  assign _zz__zz_stateReg_211 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_213 = ({1'd0,_zz_stateReg_212} <<< 1'd1);
  assign _zz__zz_stateReg_215 = ({1'd0,_zz_stateReg_214} <<< 1'd1);
  assign _zz__zz_stateReg_216 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_218 = ({1'd0,_zz_stateReg_217} <<< 1'd1);
  assign _zz__zz_stateReg_219 = ({1'd0,_zz_stateReg_79} <<< 1'd1);
  assign _zz__zz_stateReg_220 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_222 = ({1'd0,_zz_stateReg_221} <<< 1'd1);
  assign _zz__zz_stateReg_224 = ({1'd0,_zz_stateReg_223} <<< 1'd1);
  assign _zz__zz_stateReg_225 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_227 = ({1'd0,_zz_stateReg_226} <<< 1'd1);
  assign _zz__zz_stateReg_228 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_229 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_231 = ({1'd0,_zz_stateReg_230} <<< 1'd1);
  assign _zz__zz_stateReg_233 = ({1'd0,_zz_stateReg_232} <<< 1'd1);
  assign _zz__zz_stateReg_234 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_235 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_237 = ({1'd0,_zz_stateReg_236} <<< 1'd1);
  assign _zz__zz_stateReg_239 = ({1'd0,_zz_stateReg_238} <<< 1'd1);
  assign _zz__zz_stateReg_240 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_242 = ({1'd0,_zz_stateReg_241} <<< 1'd1);
  assign _zz__zz_stateReg_243 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_245 = ({1'd0,_zz_stateReg_244} <<< 1'd1);
  assign _zz__zz_stateReg_247 = ({1'd0,_zz_stateReg_246} <<< 1'd1);
  assign _zz__zz_stateReg_248 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_250 = ({1'd0,_zz_stateReg_249} <<< 1'd1);
  assign _zz__zz_stateReg_252 = ({1'd0,_zz_stateReg_251} <<< 1'd1);
  assign _zz__zz_stateReg_253 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_255 = ({1'd0,_zz_stateReg_254} <<< 1'd1);
  assign _zz__zz_stateReg_257 = ({1'd0,_zz_stateReg_256} <<< 1'd1);
  assign _zz__zz_stateReg_258 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_260 = ({1'd0,_zz_stateReg_259} <<< 1'd1);
  assign _zz__zz_stateReg_261 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_262 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_264 = ({1'd0,_zz_stateReg_263} <<< 1'd1);
  assign _zz__zz_stateReg_266 = ({1'd0,_zz_stateReg_265} <<< 1'd1);
  assign _zz__zz_stateReg_267 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_268 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_270 = ({1'd0,_zz_stateReg_269} <<< 1'd1);
  assign _zz__zz_stateReg_272 = ({1'd0,_zz_stateReg_271} <<< 1'd1);
  assign _zz__zz_stateReg_273 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_275 = ({1'd0,_zz_stateReg_274} <<< 1'd1);
  assign _zz__zz_stateReg_276 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_278 = ({1'd0,_zz_stateReg_277} <<< 1'd1);
  assign _zz__zz_stateReg_280 = ({1'd0,_zz_stateReg_279} <<< 1'd1);
  assign _zz__zz_stateReg_281 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_283 = ({1'd0,_zz_stateReg_282} <<< 1'd1);
  assign _zz__zz_stateReg_284 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_286 = ({1'd0,_zz_stateReg_285} <<< 1'd1);
  assign _zz__zz_stateReg_288 = ({1'd0,_zz_stateReg_287} <<< 1'd1);
  assign _zz__zz_stateReg_289 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_291 = ({1'd0,_zz_stateReg_290} <<< 1'd1);
  assign _zz__zz_stateReg_293 = ({1'd0,_zz_stateReg_292} <<< 1'd1);
  assign _zz__zz_stateReg_294 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_296 = ({1'd0,_zz_stateReg_295} <<< 1'd1);
  assign _zz__zz_stateReg_297 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_298 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_300 = ({1'd0,_zz_stateReg_299} <<< 1'd1);
  assign _zz__zz_stateReg_302 = ({1'd0,_zz_stateReg_301} <<< 1'd1);
  assign _zz__zz_stateReg_303 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_304 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_306 = ({1'd0,_zz_stateReg_305} <<< 1'd1);
  assign _zz__zz_stateReg_308 = ({1'd0,_zz_stateReg_307} <<< 1'd1);
  assign _zz__zz_stateReg_309 = ({1'd0,_zz_stateReg_80} <<< 1'd1);
  assign _zz__zz_stateReg_310 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_312 = ({1'd0,_zz_stateReg_311} <<< 1'd1);
  assign _zz__zz_stateReg_314 = ({1'd0,_zz_stateReg_313} <<< 1'd1);
  assign _zz__zz_stateReg_315 = ({1'd0,_zz_stateReg_81} <<< 1'd1);
  assign _zz__zz_stateReg_317 = ({1'd0,_zz_stateReg_316} <<< 1'd1);
  assign _zz__zz_stateReg_318 = ({1'd0,_zz_stateReg_82} <<< 1'd1);
  assign _zz__zz_stateReg_320 = ({1'd0,_zz_stateReg_319} <<< 1'd1);
  assign _zz__zz_stateReg_322 = ({1'd0,_zz_stateReg_321} <<< 1'd1);
  assign _zz__zz_stateReg_323 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_325 = ({1'd0,_zz_stateReg_324} <<< 1'd1);
  assign _zz__zz_stateReg_327 = ({1'd0,_zz_stateReg_326} <<< 1'd1);
  assign _zz__zz_stateReg_328 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_330 = ({1'd0,_zz_stateReg_329} <<< 1'd1);
  assign _zz__zz_stateReg_331 = ({1'd0,_zz_stateReg_83} <<< 1'd1);
  assign _zz__zz_stateReg_332 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_334 = ({1'd0,_zz_stateReg_333} <<< 1'd1);
  assign _zz__zz_stateReg_336 = ({1'd0,_zz_stateReg_335} <<< 1'd1);
  assign _zz__zz_stateReg_337 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_339 = ({1'd0,_zz_stateReg_338} <<< 1'd1);
  assign _zz__zz_stateReg_340 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_341 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_343 = ({1'd0,_zz_stateReg_342} <<< 1'd1);
  assign _zz__zz_stateReg_345 = ({1'd0,_zz_stateReg_344} <<< 1'd1);
  assign _zz__zz_stateReg_346 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_347 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_349 = ({1'd0,_zz_stateReg_348} <<< 1'd1);
  assign _zz__zz_stateReg_351 = ({1'd0,_zz_stateReg_350} <<< 1'd1);
  assign _zz__zz_stateReg_352 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_354 = ({1'd0,_zz_stateReg_353} <<< 1'd1);
  assign _zz__zz_stateReg_355 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_357 = ({1'd0,_zz_stateReg_356} <<< 1'd1);
  assign _zz__zz_stateReg_359 = ({1'd0,_zz_stateReg_358} <<< 1'd1);
  assign _zz__zz_stateReg_360 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_362 = ({1'd0,_zz_stateReg_361} <<< 1'd1);
  assign _zz__zz_stateReg_364 = ({1'd0,_zz_stateReg_363} <<< 1'd1);
  assign _zz__zz_stateReg_365 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_367 = ({1'd0,_zz_stateReg_366} <<< 1'd1);
  assign _zz__zz_stateReg_369 = ({1'd0,_zz_stateReg_368} <<< 1'd1);
  assign _zz__zz_stateReg_370 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_372 = ({1'd0,_zz_stateReg_371} <<< 1'd1);
  assign _zz__zz_stateReg_373 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_374 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_376 = ({1'd0,_zz_stateReg_375} <<< 1'd1);
  assign _zz__zz_stateReg_378 = ({1'd0,_zz_stateReg_377} <<< 1'd1);
  assign _zz__zz_stateReg_379 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_380 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_382 = ({1'd0,_zz_stateReg_381} <<< 1'd1);
  assign _zz__zz_stateReg_384 = ({1'd0,_zz_stateReg_383} <<< 1'd1);
  assign _zz__zz_stateReg_385 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_387 = ({1'd0,_zz_stateReg_386} <<< 1'd1);
  assign _zz__zz_stateReg_388 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_390 = ({1'd0,_zz_stateReg_389} <<< 1'd1);
  assign _zz__zz_stateReg_392 = ({1'd0,_zz_stateReg_391} <<< 1'd1);
  assign _zz__zz_stateReg_393 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_395 = ({1'd0,_zz_stateReg_394} <<< 1'd1);
  assign _zz__zz_stateReg_396 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_398 = ({1'd0,_zz_stateReg_397} <<< 1'd1);
  assign _zz__zz_stateReg_400 = ({1'd0,_zz_stateReg_399} <<< 1'd1);
  assign _zz__zz_stateReg_401 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_403 = ({1'd0,_zz_stateReg_402} <<< 1'd1);
  assign _zz__zz_stateReg_405 = ({1'd0,_zz_stateReg_404} <<< 1'd1);
  assign _zz__zz_stateReg_406 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_408 = ({1'd0,_zz_stateReg_407} <<< 1'd1);
  assign _zz__zz_stateReg_409 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_410 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_412 = ({1'd0,_zz_stateReg_411} <<< 1'd1);
  assign _zz__zz_stateReg_414 = ({1'd0,_zz_stateReg_413} <<< 1'd1);
  assign _zz__zz_stateReg_415 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_416 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_418 = ({1'd0,_zz_stateReg_417} <<< 1'd1);
  assign _zz__zz_stateReg_420 = ({1'd0,_zz_stateReg_419} <<< 1'd1);
  assign _zz__zz_stateReg_421 = ({1'd0,_zz_stateReg_84} <<< 1'd1);
  assign _zz__zz_stateReg_422 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_424 = ({1'd0,_zz_stateReg_423} <<< 1'd1);
  assign _zz__zz_stateReg_426 = ({1'd0,_zz_stateReg_425} <<< 1'd1);
  assign _zz__zz_stateReg_427 = ({1'd0,_zz_stateReg_85} <<< 1'd1);
  assign _zz__zz_stateReg_429 = ({1'd0,_zz_stateReg_428} <<< 1'd1);
  assign _zz__zz_stateReg_430 = ({1'd0,_zz_stateReg_86} <<< 1'd1);
  assign _zz__zz_stateReg_432 = ({1'd0,_zz_stateReg_431} <<< 1'd1);
  assign _zz__zz_stateReg_434 = ({1'd0,_zz_stateReg_433} <<< 1'd1);
  assign _zz__zz_stateReg_435 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_437 = ({1'd0,_zz_stateReg_436} <<< 1'd1);
  assign _zz__zz_stateReg_439 = ({1'd0,_zz_stateReg_438} <<< 1'd1);
  assign _zz__zz_stateReg_440 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_442 = ({1'd0,_zz_stateReg_441} <<< 1'd1);
  assign _zz__zz_stateReg_443 = ({1'd0,_zz_stateReg_87} <<< 1'd1);
  assign _zz__zz_stateReg_444 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_446 = ({1'd0,_zz_stateReg_445} <<< 1'd1);
  assign _zz__zz_stateReg_448 = ({1'd0,_zz_stateReg_447} <<< 1'd1);
  assign _zz__zz_stateReg_449 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_451 = ({1'd0,_zz_stateReg_450} <<< 1'd1);
  assign _zz__zz_stateReg_452 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_453 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_455 = ({1'd0,_zz_stateReg_454} <<< 1'd1);
  assign _zz__zz_stateReg_457 = ({1'd0,_zz_stateReg_456} <<< 1'd1);
  assign _zz__zz_stateReg_458 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_459 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_461 = ({1'd0,_zz_stateReg_460} <<< 1'd1);
  assign _zz__zz_stateReg_463 = ({1'd0,_zz_stateReg_462} <<< 1'd1);
  assign _zz__zz_stateReg_464 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_466 = ({1'd0,_zz_stateReg_465} <<< 1'd1);
  assign _zz__zz_stateReg_467 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_469 = ({1'd0,_zz_stateReg_468} <<< 1'd1);
  assign _zz__zz_stateReg_471 = ({1'd0,_zz_stateReg_470} <<< 1'd1);
  assign _zz__zz_stateReg_472 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_474 = ({1'd0,_zz_stateReg_473} <<< 1'd1);
  assign _zz__zz_stateReg_476 = ({1'd0,_zz_stateReg_475} <<< 1'd1);
  assign _zz__zz_stateReg_477 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_479 = ({1'd0,_zz_stateReg_478} <<< 1'd1);
  assign _zz__zz_stateReg_481 = ({1'd0,_zz_stateReg_480} <<< 1'd1);
  assign _zz__zz_stateReg_482 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_484 = ({1'd0,_zz_stateReg_483} <<< 1'd1);
  assign _zz__zz_stateReg_485 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_486 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_488 = ({1'd0,_zz_stateReg_487} <<< 1'd1);
  assign _zz__zz_stateReg_490 = ({1'd0,_zz_stateReg_489} <<< 1'd1);
  assign _zz__zz_stateReg_491 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_492 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_494 = ({1'd0,_zz_stateReg_493} <<< 1'd1);
  assign _zz__zz_stateReg_496 = ({1'd0,_zz_stateReg_495} <<< 1'd1);
  assign _zz__zz_stateReg_497 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_499 = ({1'd0,_zz_stateReg_498} <<< 1'd1);
  assign _zz__zz_stateReg_500 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_502 = ({1'd0,_zz_stateReg_501} <<< 1'd1);
  assign _zz__zz_stateReg_504 = ({1'd0,_zz_stateReg_503} <<< 1'd1);
  assign _zz__zz_stateReg_505 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_507 = ({1'd0,_zz_stateReg_506} <<< 1'd1);
  assign _zz__zz_stateReg_508 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_510 = ({1'd0,_zz_stateReg_509} <<< 1'd1);
  assign _zz__zz_stateReg_512 = ({1'd0,_zz_stateReg_511} <<< 1'd1);
  assign _zz__zz_stateReg_513 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_515 = ({1'd0,_zz_stateReg_514} <<< 1'd1);
  assign _zz__zz_stateReg_517 = ({1'd0,_zz_stateReg_516} <<< 1'd1);
  assign _zz__zz_stateReg_518 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_520 = ({1'd0,_zz_stateReg_519} <<< 1'd1);
  assign _zz__zz_stateReg_521 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_522 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_524 = ({1'd0,_zz_stateReg_523} <<< 1'd1);
  assign _zz__zz_stateReg_526 = ({1'd0,_zz_stateReg_525} <<< 1'd1);
  assign _zz__zz_stateReg_527 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_528 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_530 = ({1'd0,_zz_stateReg_529} <<< 1'd1);
  assign _zz__zz_stateReg_532 = ({1'd0,_zz_stateReg_531} <<< 1'd1);
  assign _zz__zz_stateReg_533 = ({1'd0,_zz_stateReg_88} <<< 1'd1);
  assign _zz__zz_stateReg_534 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_536 = ({1'd0,_zz_stateReg_535} <<< 1'd1);
  assign _zz__zz_stateReg_538 = ({1'd0,_zz_stateReg_537} <<< 1'd1);
  assign _zz__zz_stateReg_539 = ({1'd0,_zz_stateReg_89} <<< 1'd1);
  assign _zz__zz_stateReg_541 = ({1'd0,_zz_stateReg_540} <<< 1'd1);
  assign _zz__zz_stateReg_542 = ({1'd0,_zz_stateReg_90} <<< 1'd1);
  assign _zz__zz_stateReg_544 = ({1'd0,_zz_stateReg_543} <<< 1'd1);
  assign _zz__zz_stateReg_546 = ({1'd0,_zz_stateReg_545} <<< 1'd1);
  assign _zz__zz_stateReg_547 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_549 = ({1'd0,_zz_stateReg_548} <<< 1'd1);
  assign _zz__zz_stateReg_551 = ({1'd0,_zz_stateReg_550} <<< 1'd1);
  assign _zz__zz_stateReg_552 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_554 = ({1'd0,_zz_stateReg_553} <<< 1'd1);
  assign _zz__zz_stateReg_555 = ({1'd0,_zz_stateReg_91} <<< 1'd1);
  assign _zz__zz_stateReg_4_1 = stateReg[127 : 120];
  assign _zz__zz_stateReg_8_1 = stateReg[95 : 88];
  assign _zz__zz_stateReg_12_1 = stateReg[63 : 56];
  assign _zz__zz_stateReg_16_1 = stateReg[31 : 24];
  assign _zz__zz_stateReg_5_1 = stateReg[87 : 80];
  assign _zz__zz_stateReg_9_1 = stateReg[55 : 48];
  assign _zz__zz_stateReg_13_1 = stateReg[23 : 16];
  assign _zz__zz_stateReg_17_1 = stateReg[119 : 112];
  assign _zz__zz_stateReg_6_1 = stateReg[47 : 40];
  assign _zz__zz_stateReg_10_1 = stateReg[15 : 8];
  assign _zz__zz_stateReg_14_1 = stateReg[111 : 104];
  assign _zz__zz_stateReg_18_1 = stateReg[79 : 72];
  assign _zz__zz_stateReg_7_1 = stateReg[7 : 0];
  assign _zz__zz_stateReg_11_1 = stateReg[103 : 96];
  assign _zz__zz_stateReg_15_1 = stateReg[71 : 64];
  assign _zz__zz_stateReg_19_1 = stateReg[39 : 32];
  assign _zz__zz_roundKeyReg_0_2_1 = _zz_roundKeyReg_0_1[31 : 24];
  assign _zz__zz_roundKeyReg_0_2_3 = _zz_roundKeyReg_0_1[23 : 16];
  assign _zz__zz_roundKeyReg_0_2_5 = _zz_roundKeyReg_0_1[15 : 8];
  assign _zz__zz_roundKeyReg_0_2_7 = _zz_roundKeyReg_0_1[7 : 0];
  assign _zz__zz_stateReg_71_1 = _zz_stateReg_70[31 : 24];
  assign _zz__zz_stateReg_71_3 = _zz_stateReg_70[23 : 16];
  assign _zz__zz_stateReg_71_5 = _zz_stateReg_70[15 : 8];
  assign _zz__zz_stateReg_71_7 = _zz_stateReg_70[7 : 0];
  assign _zz__zz_roundKeyReg_0_4_1 = _zz_roundKeyReg_0_3[31 : 24];
  assign _zz__zz_roundKeyReg_0_4_3 = _zz_roundKeyReg_0_3[23 : 16];
  assign _zz__zz_roundKeyReg_0_4_5 = _zz_roundKeyReg_0_3[15 : 8];
  assign _zz__zz_roundKeyReg_0_4_7 = _zz_roundKeyReg_0_3[7 : 0];
  assign _zz__zz_stateReg_75_3 = stateReg[127 : 120];
  assign _zz__zz_stateReg_75_5 = stateReg[23 : 16];
  assign _zz__zz_stateReg_75_7 = stateReg[47 : 40];
  assign _zz__zz_stateReg_75_9 = stateReg[71 : 64];
  assign _zz__zz_stateReg_75_12 = stateReg[95 : 88];
  assign _zz__zz_stateReg_75_14 = stateReg[119 : 112];
  assign _zz__zz_stateReg_75_16 = stateReg[15 : 8];
  assign _zz__zz_stateReg_75_18 = stateReg[39 : 32];
  assign _zz__zz_stateReg_75_20 = stateReg[63 : 56];
  assign _zz__zz_stateReg_75_22 = stateReg[87 : 80];
  assign _zz__zz_stateReg_75_25 = stateReg[111 : 104];
  assign _zz__zz_stateReg_75_27 = stateReg[7 : 0];
  assign _zz__zz_stateReg_75_29 = stateReg[31 : 24];
  assign _zz__zz_stateReg_75_31 = stateReg[55 : 48];
  assign _zz__zz_stateReg_75_33 = stateReg[79 : 72];
  assign _zz__zz_stateReg_75_35 = stateReg[103 : 96];
  assign _zz_stateReg_556 = {{{{{_zz_stateReg_557,_zz_stateReg_563},_zz_stateReg_564},(_zz_stateReg_565 ^ _zz_stateReg_566)},(_zz_stateReg_567 ^ _zz_stateReg_2[31 : 24])},(io_dataIn[55 : 48] ^ _zz_stateReg_2[23 : 16])};
  assign _zz_stateReg_568 = (io_dataIn[47 : 40] ^ _zz_stateReg_2[15 : 8]);
  assign _zz_stateReg_569 = (io_dataIn[39 : 32] ^ _zz_stateReg_2[7 : 0]);
  assign _zz_stateReg_570 = io_dataIn[31 : 24];
  assign _zz_stateReg_571 = _zz_stateReg_3[31 : 24];
  assign _zz_stateReg_572 = io_dataIn[23 : 16];
  assign _zz_stateReg_557 = {{{{_zz_stateReg_558,_zz_stateReg_559},(_zz_stateReg_560 ^ _zz_stateReg_561)},(_zz_stateReg_562 ^ _zz_stateReg[7 : 0])},(io_dataIn[95 : 88] ^ _zz_stateReg_1[31 : 24])};
  assign _zz_stateReg_563 = (io_dataIn[87 : 80] ^ _zz_stateReg_1[23 : 16]);
  assign _zz_stateReg_564 = (io_dataIn[79 : 72] ^ _zz_stateReg_1[15 : 8]);
  assign _zz_stateReg_565 = io_dataIn[71 : 64];
  assign _zz_stateReg_566 = _zz_stateReg_1[7 : 0];
  assign _zz_stateReg_567 = io_dataIn[63 : 56];
  assign _zz_stateReg_558 = (io_dataIn[127 : 120] ^ _zz_stateReg[31 : 24]);
  assign _zz_stateReg_559 = (io_dataIn[119 : 112] ^ _zz_stateReg[23 : 16]);
  assign _zz_stateReg_560 = io_dataIn[111 : 104];
  assign _zz_stateReg_561 = _zz_stateReg[15 : 8];
  assign _zz_stateReg_562 = io_dataIn[103 : 96];
  assign _zz__zz_stateReg_68 = {{{{_zz_stateReg_20,_zz_stateReg_21},_zz_stateReg_22},_zz_stateReg_23},_zz_stateReg_24};
  assign _zz__zz_stateReg_68_1 = _zz_stateReg_25;
  assign _zz__zz_stateReg_69 = {{{{{{_zz_roundKeyReg_0_2[31 : 24],_zz_roundKeyReg_0_2[23 : 16]},_zz_roundKeyReg_0_2[15 : 8]},_zz_roundKeyReg_0_2[7 : 0]},_zz_roundKeyReg_1[31 : 24]},_zz_roundKeyReg_1[23 : 16]},_zz_roundKeyReg_1[15 : 8]};
  assign _zz__zz_stateReg_69_1 = _zz_roundKeyReg_1[7 : 0];
  assign _zz__zz_stateReg_69_2 = _zz_roundKeyReg_2[31 : 24];
  assign _zz_stateReg_573 = {{{{{{_zz_stateReg_71[31 : 24],_zz_stateReg_71[23 : 16]},_zz_stateReg_71[15 : 8]},_zz_stateReg_71[7 : 0]},_zz_stateReg_72[31 : 24]},_zz_stateReg_72[23 : 16]},_zz_stateReg_72[15 : 8]};
  assign _zz_stateReg_574 = _zz_stateReg_72[7 : 0];
  assign _zz_stateReg_575 = _zz_stateReg_73[31 : 24];
  assign _zz__zz_stateReg_75 = {{{{{{_zz__zz_stateReg_75_1,_zz__zz_stateReg_75_10},_zz__zz_stateReg_75_13},_zz__zz_stateReg_75_15},_zz__zz_stateReg_75_17},_zz__zz_stateReg_75_19},_zz__zz_stateReg_75_21};
  assign _zz__zz_stateReg_75_23 = _zz__zz_stateReg_75_24;
  assign _zz__zz_stateReg_75_36 = {{{{{{_zz__zz_stateReg_75_37,_zz__zz_stateReg_75_38},_zz__zz_stateReg_75_39},_zz_roundKeyReg_1_1[15 : 8]},_zz_roundKeyReg_1_1[7 : 0]},_zz_roundKeyReg_2_1[31 : 24]},_zz_roundKeyReg_2_1[23 : 16]};
  assign _zz__zz_stateReg_75_40 = _zz_roundKeyReg_2_1[15 : 8];
  assign _zz__zz_stateReg_75_41 = _zz_roundKeyReg_2_1[7 : 0];
  assign _zz__zz_stateReg_75_1 = {{{_zz__zz_stateReg_75_2,_zz__zz_stateReg_75_4},_zz__zz_stateReg_75_6},_zz__zz_stateReg_75_8};
  assign _zz__zz_stateReg_75_10 = _zz__zz_stateReg_75_11;
  assign _zz__zz_stateReg_75_37 = {{{_zz_roundKeyReg_0_4[31 : 24],_zz_roundKeyReg_0_4[23 : 16]},_zz_roundKeyReg_0_4[15 : 8]},_zz_roundKeyReg_0_4[7 : 0]};
  assign _zz__zz_stateReg_75_38 = _zz_roundKeyReg_1_1[31 : 24];
  assign _zz__zz_stateReg_75_39 = _zz_roundKeyReg_1_1[23 : 16];
  assign _zz__zz_stateReg_92 = (_zz_stateReg_111[7] ? (_zz_stateReg_112 ^ 8'h1b) : _zz_stateReg_112);
  assign _zz__zz_stateReg_92_1 = (_zz_stateReg_114[7] ? (_zz_stateReg_115 ^ 8'h1b) : _zz_stateReg_115);
  assign _zz__zz_stateReg_92_2 = _zz_stateReg_76[7];
  assign _zz__zz_stateReg_92_3 = (_zz_stateReg_116 ^ 8'h1b);
  assign _zz__zz_stateReg_92_4 = (_zz_stateReg_120[7] ? (_zz_stateReg_121 ^ 8'h1b) : _zz_stateReg_121);
  assign _zz__zz_stateReg_92_5 = (_zz_stateReg_77[7] ? (_zz_stateReg_122 ^ 8'h1b) : _zz_stateReg_122);
  assign _zz__zz_stateReg_92_6 = _zz_stateReg_126[7];
  assign _zz__zz_stateReg_92_7 = (_zz_stateReg_127 ^ 8'h1b);
  assign _zz__zz_stateReg_92_8 = _zz_stateReg_129[7];
  assign _zz__zz_stateReg_92_9 = (_zz_stateReg_130 ^ 8'h1b);
  assign _zz__zz_stateReg_93 = _zz_stateReg_139[7];
  assign _zz__zz_stateReg_93_1 = (_zz_stateReg_140 ^ 8'h1b);
  assign _zz__zz_stateReg_93_2 = (_zz_stateReg_144[7] ? (_zz_stateReg_145 ^ 8'h1b) : _zz_stateReg_145);
  assign _zz__zz_stateReg_93_3 = (_zz_stateReg_147[7] ? (_zz_stateReg_148 ^ 8'h1b) : _zz_stateReg_148);
  assign _zz__zz_stateReg_93_4 = _zz_stateReg_77[7];
  assign _zz__zz_stateReg_93_5 = (_zz_stateReg_149 ^ 8'h1b);
  assign _zz__zz_stateReg_93_6 = _zz_stateReg_153[7];
  assign _zz__zz_stateReg_93_7 = (_zz_stateReg_154 ^ 8'h1b);
  assign _zz__zz_stateReg_93_8 = _zz_stateReg_78[7];
  assign _zz__zz_stateReg_93_9 = (_zz_stateReg_155 ^ 8'h1b);
  assign _zz__zz_stateReg_93_10 = 8'h1b;
  assign _zz__zz_stateReg_93_11 = 8'h1b;
  assign _zz__zz_stateReg_94 = (_zz_stateReg_167[7] ? (_zz_stateReg_168 ^ 8'h1b) : _zz_stateReg_168);
  assign _zz__zz_stateReg_94_1 = (_zz_stateReg_170[7] ? (_zz_stateReg_171 ^ 8'h1b) : _zz_stateReg_171);
  assign _zz__zz_stateReg_94_2 = _zz_stateReg_175[7];
  assign _zz__zz_stateReg_94_3 = (_zz_stateReg_176 ^ 8'h1b);
  assign _zz__zz_stateReg_94_4 = _zz_stateReg_180[7];
  assign _zz__zz_stateReg_94_5 = (_zz_stateReg_181 ^ 8'h1b);
  assign _zz__zz_stateReg_94_6 = _zz_stateReg_183[7];
  assign _zz__zz_stateReg_94_7 = (_zz_stateReg_184 ^ 8'h1b);
  assign _zz__zz_stateReg_94_8 = 8'h1b;
  assign _zz__zz_stateReg_94_9 = 8'h1b;
  assign _zz__zz_stateReg_94_10 = 8'h1b;
  assign _zz__zz_stateReg_95 = (_zz_stateReg_195[7] ? (_zz_stateReg_196 ^ 8'h1b) : _zz_stateReg_196);
  assign _zz__zz_stateReg_95_1 = (_zz_stateReg_76[7] ? (_zz_stateReg_197 ^ 8'h1b) : _zz_stateReg_197);
  assign _zz__zz_stateReg_95_2 = (_zz_stateReg_201[7] ? (_zz_stateReg_202 ^ 8'h1b) : _zz_stateReg_202);
  assign _zz__zz_stateReg_95_3 = (_zz_stateReg_204[7] ? (_zz_stateReg_205 ^ 8'h1b) : _zz_stateReg_205);
  assign _zz__zz_stateReg_95_4 = 8'h1b;
  assign _zz__zz_stateReg_95_5 = 8'h1b;
  assign _zz__zz_stateReg_95_6 = 8'h1b;
  assign _zz__zz_stateReg_96 = (_zz_stateReg_223[7] ? (_zz_stateReg_224 ^ 8'h1b) : _zz_stateReg_224);
  assign _zz__zz_stateReg_96_1 = (_zz_stateReg_226[7] ? (_zz_stateReg_227 ^ 8'h1b) : _zz_stateReg_227);
  assign _zz__zz_stateReg_96_2 = _zz_stateReg_80[7];
  assign _zz__zz_stateReg_96_3 = (_zz_stateReg_228 ^ 8'h1b);
  assign _zz__zz_stateReg_96_4 = (_zz_stateReg_232[7] ? (_zz_stateReg_233 ^ 8'h1b) : _zz_stateReg_233);
  assign _zz__zz_stateReg_96_5 = (_zz_stateReg_81[7] ? (_zz_stateReg_234 ^ 8'h1b) : _zz_stateReg_234);
  assign _zz__zz_stateReg_96_6 = _zz_stateReg_238[7];
  assign _zz__zz_stateReg_96_7 = (_zz_stateReg_239 ^ 8'h1b);
  assign _zz__zz_stateReg_96_8 = _zz_stateReg_241[7];
  assign _zz__zz_stateReg_96_9 = (_zz_stateReg_242 ^ 8'h1b);
  assign _zz__zz_stateReg_97 = _zz_stateReg_251[7];
  assign _zz__zz_stateReg_97_1 = (_zz_stateReg_252 ^ 8'h1b);
  assign _zz__zz_stateReg_97_2 = (_zz_stateReg_256[7] ? (_zz_stateReg_257 ^ 8'h1b) : _zz_stateReg_257);
  assign _zz__zz_stateReg_97_3 = (_zz_stateReg_259[7] ? (_zz_stateReg_260 ^ 8'h1b) : _zz_stateReg_260);
  assign _zz__zz_stateReg_97_4 = _zz_stateReg_81[7];
  assign _zz__zz_stateReg_97_5 = (_zz_stateReg_261 ^ 8'h1b);
  assign _zz__zz_stateReg_97_6 = _zz_stateReg_265[7];
  assign _zz__zz_stateReg_97_7 = (_zz_stateReg_266 ^ 8'h1b);
  assign _zz__zz_stateReg_97_8 = _zz_stateReg_82[7];
  assign _zz__zz_stateReg_97_9 = (_zz_stateReg_267 ^ 8'h1b);
  assign _zz__zz_stateReg_97_10 = 8'h1b;
  assign _zz__zz_stateReg_97_11 = 8'h1b;
  assign _zz__zz_stateReg_98 = (_zz_stateReg_279[7] ? (_zz_stateReg_280 ^ 8'h1b) : _zz_stateReg_280);
  assign _zz__zz_stateReg_98_1 = (_zz_stateReg_282[7] ? (_zz_stateReg_283 ^ 8'h1b) : _zz_stateReg_283);
  assign _zz__zz_stateReg_98_2 = _zz_stateReg_287[7];
  assign _zz__zz_stateReg_98_3 = (_zz_stateReg_288 ^ 8'h1b);
  assign _zz__zz_stateReg_98_4 = _zz_stateReg_292[7];
  assign _zz__zz_stateReg_98_5 = (_zz_stateReg_293 ^ 8'h1b);
  assign _zz__zz_stateReg_98_6 = _zz_stateReg_295[7];
  assign _zz__zz_stateReg_98_7 = (_zz_stateReg_296 ^ 8'h1b);
  assign _zz__zz_stateReg_98_8 = 8'h1b;
  assign _zz__zz_stateReg_98_9 = 8'h1b;
  assign _zz__zz_stateReg_98_10 = 8'h1b;
  assign _zz__zz_stateReg_99 = (_zz_stateReg_307[7] ? (_zz_stateReg_308 ^ 8'h1b) : _zz_stateReg_308);
  assign _zz__zz_stateReg_99_1 = (_zz_stateReg_80[7] ? (_zz_stateReg_309 ^ 8'h1b) : _zz_stateReg_309);
  assign _zz__zz_stateReg_99_2 = (_zz_stateReg_313[7] ? (_zz_stateReg_314 ^ 8'h1b) : _zz_stateReg_314);
  assign _zz__zz_stateReg_99_3 = (_zz_stateReg_316[7] ? (_zz_stateReg_317 ^ 8'h1b) : _zz_stateReg_317);
  assign _zz__zz_stateReg_99_4 = 8'h1b;
  assign _zz__zz_stateReg_99_5 = 8'h1b;
  assign _zz__zz_stateReg_99_6 = 8'h1b;
  assign _zz__zz_stateReg_100 = (_zz_stateReg_335[7] ? (_zz_stateReg_336 ^ 8'h1b) : _zz_stateReg_336);
  assign _zz__zz_stateReg_100_1 = (_zz_stateReg_338[7] ? (_zz_stateReg_339 ^ 8'h1b) : _zz_stateReg_339);
  assign _zz__zz_stateReg_100_2 = _zz_stateReg_84[7];
  assign _zz__zz_stateReg_100_3 = (_zz_stateReg_340 ^ 8'h1b);
  assign _zz__zz_stateReg_100_4 = (_zz_stateReg_344[7] ? (_zz_stateReg_345 ^ 8'h1b) : _zz_stateReg_345);
  assign _zz__zz_stateReg_100_5 = (_zz_stateReg_85[7] ? (_zz_stateReg_346 ^ 8'h1b) : _zz_stateReg_346);
  assign _zz__zz_stateReg_100_6 = _zz_stateReg_350[7];
  assign _zz__zz_stateReg_100_7 = (_zz_stateReg_351 ^ 8'h1b);
  assign _zz__zz_stateReg_100_8 = _zz_stateReg_353[7];
  assign _zz__zz_stateReg_100_9 = (_zz_stateReg_354 ^ 8'h1b);
  assign _zz__zz_stateReg_101 = _zz_stateReg_363[7];
  assign _zz__zz_stateReg_101_1 = (_zz_stateReg_364 ^ 8'h1b);
  assign _zz__zz_stateReg_101_2 = (_zz_stateReg_368[7] ? (_zz_stateReg_369 ^ 8'h1b) : _zz_stateReg_369);
  assign _zz__zz_stateReg_101_3 = (_zz_stateReg_371[7] ? (_zz_stateReg_372 ^ 8'h1b) : _zz_stateReg_372);
  assign _zz__zz_stateReg_101_4 = _zz_stateReg_85[7];
  assign _zz__zz_stateReg_101_5 = (_zz_stateReg_373 ^ 8'h1b);
  assign _zz__zz_stateReg_101_6 = _zz_stateReg_377[7];
  assign _zz__zz_stateReg_101_7 = (_zz_stateReg_378 ^ 8'h1b);
  assign _zz__zz_stateReg_101_8 = _zz_stateReg_86[7];
  assign _zz__zz_stateReg_101_9 = (_zz_stateReg_379 ^ 8'h1b);
  assign _zz__zz_stateReg_101_10 = 8'h1b;
  assign _zz__zz_stateReg_101_11 = 8'h1b;
  assign _zz__zz_stateReg_102 = (_zz_stateReg_391[7] ? (_zz_stateReg_392 ^ 8'h1b) : _zz_stateReg_392);
  assign _zz__zz_stateReg_102_1 = (_zz_stateReg_394[7] ? (_zz_stateReg_395 ^ 8'h1b) : _zz_stateReg_395);
  assign _zz__zz_stateReg_102_2 = _zz_stateReg_399[7];
  assign _zz__zz_stateReg_102_3 = (_zz_stateReg_400 ^ 8'h1b);
  assign _zz__zz_stateReg_102_4 = _zz_stateReg_404[7];
  assign _zz__zz_stateReg_102_5 = (_zz_stateReg_405 ^ 8'h1b);
  assign _zz__zz_stateReg_102_6 = _zz_stateReg_407[7];
  assign _zz__zz_stateReg_102_7 = (_zz_stateReg_408 ^ 8'h1b);
  assign _zz__zz_stateReg_102_8 = 8'h1b;
  assign _zz__zz_stateReg_102_9 = 8'h1b;
  assign _zz__zz_stateReg_102_10 = 8'h1b;
  assign _zz__zz_stateReg_103 = (_zz_stateReg_419[7] ? (_zz_stateReg_420 ^ 8'h1b) : _zz_stateReg_420);
  assign _zz__zz_stateReg_103_1 = (_zz_stateReg_84[7] ? (_zz_stateReg_421 ^ 8'h1b) : _zz_stateReg_421);
  assign _zz__zz_stateReg_103_2 = (_zz_stateReg_425[7] ? (_zz_stateReg_426 ^ 8'h1b) : _zz_stateReg_426);
  assign _zz__zz_stateReg_103_3 = (_zz_stateReg_428[7] ? (_zz_stateReg_429 ^ 8'h1b) : _zz_stateReg_429);
  assign _zz__zz_stateReg_103_4 = 8'h1b;
  assign _zz__zz_stateReg_103_5 = 8'h1b;
  assign _zz__zz_stateReg_103_6 = 8'h1b;
  assign _zz__zz_stateReg_104 = (_zz_stateReg_447[7] ? (_zz_stateReg_448 ^ 8'h1b) : _zz_stateReg_448);
  assign _zz__zz_stateReg_104_1 = (_zz_stateReg_450[7] ? (_zz_stateReg_451 ^ 8'h1b) : _zz_stateReg_451);
  assign _zz__zz_stateReg_104_2 = _zz_stateReg_88[7];
  assign _zz__zz_stateReg_104_3 = (_zz_stateReg_452 ^ 8'h1b);
  assign _zz__zz_stateReg_104_4 = (_zz_stateReg_456[7] ? (_zz_stateReg_457 ^ 8'h1b) : _zz_stateReg_457);
  assign _zz__zz_stateReg_104_5 = (_zz_stateReg_89[7] ? (_zz_stateReg_458 ^ 8'h1b) : _zz_stateReg_458);
  assign _zz__zz_stateReg_104_6 = _zz_stateReg_462[7];
  assign _zz__zz_stateReg_104_7 = (_zz_stateReg_463 ^ 8'h1b);
  assign _zz__zz_stateReg_104_8 = _zz_stateReg_465[7];
  assign _zz__zz_stateReg_104_9 = (_zz_stateReg_466 ^ 8'h1b);
  assign _zz__zz_stateReg_105 = _zz_stateReg_475[7];
  assign _zz__zz_stateReg_105_1 = (_zz_stateReg_476 ^ 8'h1b);
  assign _zz__zz_stateReg_105_2 = (_zz_stateReg_480[7] ? (_zz_stateReg_481 ^ 8'h1b) : _zz_stateReg_481);
  assign _zz__zz_stateReg_105_3 = (_zz_stateReg_483[7] ? (_zz_stateReg_484 ^ 8'h1b) : _zz_stateReg_484);
  assign _zz__zz_stateReg_105_4 = _zz_stateReg_89[7];
  assign _zz__zz_stateReg_105_5 = (_zz_stateReg_485 ^ 8'h1b);
  assign _zz__zz_stateReg_105_6 = _zz_stateReg_489[7];
  assign _zz__zz_stateReg_105_7 = (_zz_stateReg_490 ^ 8'h1b);
  assign _zz__zz_stateReg_105_8 = _zz_stateReg_90[7];
  assign _zz__zz_stateReg_105_9 = (_zz_stateReg_491 ^ 8'h1b);
  assign _zz__zz_stateReg_105_10 = 8'h1b;
  assign _zz__zz_stateReg_105_11 = 8'h1b;
  assign _zz__zz_stateReg_106 = (_zz_stateReg_503[7] ? (_zz_stateReg_504 ^ 8'h1b) : _zz_stateReg_504);
  assign _zz__zz_stateReg_106_1 = (_zz_stateReg_506[7] ? (_zz_stateReg_507 ^ 8'h1b) : _zz_stateReg_507);
  assign _zz__zz_stateReg_106_2 = _zz_stateReg_511[7];
  assign _zz__zz_stateReg_106_3 = (_zz_stateReg_512 ^ 8'h1b);
  assign _zz__zz_stateReg_106_4 = _zz_stateReg_516[7];
  assign _zz__zz_stateReg_106_5 = (_zz_stateReg_517 ^ 8'h1b);
  assign _zz__zz_stateReg_106_6 = _zz_stateReg_519[7];
  assign _zz__zz_stateReg_106_7 = (_zz_stateReg_520 ^ 8'h1b);
  assign _zz__zz_stateReg_106_8 = 8'h1b;
  assign _zz__zz_stateReg_106_9 = 8'h1b;
  assign _zz__zz_stateReg_106_10 = 8'h1b;
  assign _zz__zz_stateReg_107 = (_zz_stateReg_531[7] ? (_zz_stateReg_532 ^ 8'h1b) : _zz_stateReg_532);
  assign _zz__zz_stateReg_107_1 = (_zz_stateReg_88[7] ? (_zz_stateReg_533 ^ 8'h1b) : _zz_stateReg_533);
  assign _zz__zz_stateReg_107_2 = (_zz_stateReg_537[7] ? (_zz_stateReg_538 ^ 8'h1b) : _zz_stateReg_538);
  assign _zz__zz_stateReg_107_3 = (_zz_stateReg_540[7] ? (_zz_stateReg_541 ^ 8'h1b) : _zz_stateReg_541);
  assign _zz__zz_stateReg_107_4 = 8'h1b;
  assign _zz__zz_stateReg_107_5 = 8'h1b;
  assign _zz__zz_stateReg_107_6 = 8'h1b;
  assign _zz_stateReg_576 = {{{{_zz_stateReg_92,_zz_stateReg_93},_zz_stateReg_94},_zz_stateReg_95},_zz_stateReg_96};
  assign _zz_stateReg_577 = _zz_stateReg_97;
  always @(*) begin
    case(_zz__zz_stateReg_4_1)
      8'b00000000 : _zz__zz_stateReg_4 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_4 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_4 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_4 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_4 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_4 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_4 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_4 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_4 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_4 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_4 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_4 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_4 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_4 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_4 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_4 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_4 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_4 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_4 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_4 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_4 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_4 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_4 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_4 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_4 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_4 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_4 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_4 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_4 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_4 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_4 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_4 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_4 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_4 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_4 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_4 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_4 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_4 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_4 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_4 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_4 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_4 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_4 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_4 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_4 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_4 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_4 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_4 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_4 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_4 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_4 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_4 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_4 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_4 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_4 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_4 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_4 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_4 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_4 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_4 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_4 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_4 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_4 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_4 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_4 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_4 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_4 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_4 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_4 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_4 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_4 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_4 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_4 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_4 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_4 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_4 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_4 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_4 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_4 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_4 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_4 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_4 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_4 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_4 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_4 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_4 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_4 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_4 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_4 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_4 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_4 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_4 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_4 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_4 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_4 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_4 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_4 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_4 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_4 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_4 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_4 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_4 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_4 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_4 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_4 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_4 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_4 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_4 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_4 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_4 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_4 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_4 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_4 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_4 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_4 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_4 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_4 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_4 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_4 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_4 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_4 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_4 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_4 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_4 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_4 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_4 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_4 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_4 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_4 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_4 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_4 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_4 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_4 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_4 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_4 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_4 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_4 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_4 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_4 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_4 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_4 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_4 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_4 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_4 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_4 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_4 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_4 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_4 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_4 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_4 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_4 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_4 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_4 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_4 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_4 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_4 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_4 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_4 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_4 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_4 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_4 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_4 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_4 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_4 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_4 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_4 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_4 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_4 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_4 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_4 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_4 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_4 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_4 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_4 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_4 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_4 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_4 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_4 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_4 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_4 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_4 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_4 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_4 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_4 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_4 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_4 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_4 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_4 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_4 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_4 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_4 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_4 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_4 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_4 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_4 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_4 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_4 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_4 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_4 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_4 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_4 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_4 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_4 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_4 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_4 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_4 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_4 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_4 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_4 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_4 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_4 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_4 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_4 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_4 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_4 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_4 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_4 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_4 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_4 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_4 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_4 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_4 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_4 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_4 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_4 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_4 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_4 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_4 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_4 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_4 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_4 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_4 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_4 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_4 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_4 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_4 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_4 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_4 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_4 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_4 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_4 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_4 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_4 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_4 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_4 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_4 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_4 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_4 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_4 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_4 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_4 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_4 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_4 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_4 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_4 = sboxRom_254;
      default : _zz__zz_stateReg_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_8_1)
      8'b00000000 : _zz__zz_stateReg_8 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_8 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_8 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_8 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_8 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_8 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_8 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_8 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_8 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_8 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_8 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_8 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_8 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_8 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_8 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_8 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_8 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_8 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_8 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_8 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_8 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_8 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_8 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_8 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_8 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_8 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_8 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_8 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_8 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_8 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_8 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_8 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_8 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_8 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_8 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_8 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_8 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_8 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_8 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_8 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_8 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_8 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_8 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_8 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_8 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_8 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_8 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_8 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_8 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_8 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_8 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_8 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_8 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_8 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_8 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_8 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_8 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_8 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_8 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_8 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_8 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_8 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_8 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_8 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_8 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_8 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_8 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_8 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_8 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_8 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_8 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_8 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_8 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_8 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_8 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_8 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_8 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_8 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_8 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_8 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_8 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_8 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_8 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_8 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_8 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_8 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_8 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_8 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_8 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_8 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_8 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_8 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_8 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_8 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_8 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_8 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_8 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_8 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_8 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_8 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_8 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_8 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_8 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_8 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_8 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_8 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_8 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_8 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_8 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_8 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_8 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_8 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_8 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_8 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_8 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_8 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_8 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_8 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_8 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_8 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_8 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_8 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_8 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_8 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_8 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_8 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_8 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_8 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_8 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_8 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_8 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_8 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_8 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_8 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_8 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_8 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_8 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_8 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_8 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_8 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_8 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_8 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_8 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_8 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_8 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_8 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_8 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_8 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_8 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_8 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_8 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_8 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_8 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_8 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_8 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_8 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_8 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_8 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_8 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_8 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_8 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_8 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_8 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_8 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_8 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_8 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_8 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_8 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_8 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_8 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_8 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_8 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_8 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_8 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_8 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_8 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_8 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_8 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_8 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_8 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_8 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_8 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_8 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_8 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_8 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_8 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_8 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_8 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_8 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_8 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_8 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_8 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_8 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_8 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_8 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_8 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_8 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_8 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_8 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_8 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_8 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_8 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_8 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_8 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_8 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_8 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_8 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_8 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_8 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_8 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_8 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_8 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_8 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_8 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_8 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_8 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_8 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_8 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_8 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_8 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_8 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_8 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_8 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_8 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_8 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_8 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_8 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_8 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_8 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_8 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_8 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_8 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_8 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_8 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_8 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_8 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_8 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_8 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_8 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_8 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_8 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_8 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_8 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_8 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_8 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_8 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_8 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_8 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_8 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_8 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_8 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_8 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_8 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_8 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_8 = sboxRom_254;
      default : _zz__zz_stateReg_8 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_12_1)
      8'b00000000 : _zz__zz_stateReg_12 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_12 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_12 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_12 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_12 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_12 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_12 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_12 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_12 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_12 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_12 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_12 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_12 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_12 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_12 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_12 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_12 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_12 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_12 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_12 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_12 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_12 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_12 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_12 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_12 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_12 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_12 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_12 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_12 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_12 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_12 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_12 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_12 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_12 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_12 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_12 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_12 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_12 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_12 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_12 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_12 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_12 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_12 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_12 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_12 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_12 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_12 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_12 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_12 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_12 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_12 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_12 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_12 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_12 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_12 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_12 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_12 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_12 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_12 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_12 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_12 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_12 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_12 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_12 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_12 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_12 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_12 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_12 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_12 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_12 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_12 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_12 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_12 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_12 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_12 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_12 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_12 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_12 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_12 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_12 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_12 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_12 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_12 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_12 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_12 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_12 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_12 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_12 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_12 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_12 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_12 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_12 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_12 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_12 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_12 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_12 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_12 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_12 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_12 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_12 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_12 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_12 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_12 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_12 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_12 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_12 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_12 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_12 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_12 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_12 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_12 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_12 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_12 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_12 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_12 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_12 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_12 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_12 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_12 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_12 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_12 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_12 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_12 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_12 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_12 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_12 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_12 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_12 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_12 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_12 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_12 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_12 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_12 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_12 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_12 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_12 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_12 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_12 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_12 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_12 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_12 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_12 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_12 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_12 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_12 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_12 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_12 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_12 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_12 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_12 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_12 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_12 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_12 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_12 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_12 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_12 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_12 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_12 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_12 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_12 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_12 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_12 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_12 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_12 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_12 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_12 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_12 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_12 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_12 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_12 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_12 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_12 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_12 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_12 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_12 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_12 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_12 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_12 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_12 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_12 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_12 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_12 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_12 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_12 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_12 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_12 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_12 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_12 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_12 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_12 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_12 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_12 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_12 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_12 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_12 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_12 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_12 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_12 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_12 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_12 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_12 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_12 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_12 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_12 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_12 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_12 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_12 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_12 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_12 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_12 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_12 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_12 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_12 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_12 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_12 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_12 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_12 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_12 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_12 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_12 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_12 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_12 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_12 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_12 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_12 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_12 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_12 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_12 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_12 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_12 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_12 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_12 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_12 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_12 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_12 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_12 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_12 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_12 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_12 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_12 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_12 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_12 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_12 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_12 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_12 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_12 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_12 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_12 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_12 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_12 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_12 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_12 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_12 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_12 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_12 = sboxRom_254;
      default : _zz__zz_stateReg_12 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_16_1)
      8'b00000000 : _zz__zz_stateReg_16 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_16 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_16 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_16 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_16 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_16 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_16 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_16 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_16 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_16 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_16 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_16 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_16 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_16 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_16 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_16 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_16 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_16 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_16 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_16 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_16 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_16 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_16 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_16 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_16 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_16 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_16 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_16 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_16 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_16 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_16 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_16 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_16 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_16 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_16 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_16 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_16 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_16 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_16 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_16 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_16 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_16 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_16 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_16 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_16 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_16 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_16 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_16 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_16 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_16 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_16 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_16 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_16 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_16 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_16 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_16 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_16 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_16 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_16 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_16 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_16 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_16 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_16 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_16 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_16 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_16 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_16 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_16 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_16 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_16 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_16 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_16 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_16 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_16 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_16 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_16 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_16 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_16 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_16 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_16 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_16 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_16 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_16 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_16 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_16 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_16 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_16 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_16 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_16 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_16 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_16 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_16 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_16 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_16 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_16 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_16 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_16 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_16 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_16 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_16 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_16 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_16 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_16 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_16 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_16 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_16 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_16 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_16 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_16 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_16 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_16 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_16 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_16 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_16 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_16 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_16 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_16 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_16 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_16 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_16 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_16 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_16 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_16 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_16 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_16 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_16 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_16 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_16 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_16 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_16 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_16 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_16 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_16 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_16 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_16 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_16 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_16 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_16 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_16 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_16 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_16 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_16 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_16 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_16 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_16 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_16 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_16 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_16 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_16 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_16 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_16 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_16 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_16 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_16 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_16 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_16 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_16 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_16 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_16 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_16 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_16 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_16 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_16 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_16 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_16 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_16 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_16 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_16 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_16 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_16 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_16 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_16 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_16 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_16 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_16 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_16 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_16 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_16 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_16 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_16 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_16 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_16 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_16 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_16 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_16 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_16 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_16 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_16 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_16 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_16 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_16 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_16 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_16 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_16 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_16 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_16 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_16 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_16 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_16 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_16 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_16 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_16 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_16 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_16 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_16 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_16 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_16 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_16 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_16 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_16 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_16 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_16 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_16 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_16 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_16 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_16 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_16 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_16 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_16 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_16 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_16 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_16 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_16 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_16 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_16 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_16 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_16 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_16 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_16 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_16 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_16 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_16 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_16 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_16 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_16 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_16 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_16 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_16 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_16 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_16 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_16 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_16 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_16 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_16 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_16 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_16 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_16 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_16 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_16 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_16 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_16 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_16 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_16 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_16 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_16 = sboxRom_254;
      default : _zz__zz_stateReg_16 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_5_1)
      8'b00000000 : _zz__zz_stateReg_5 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_5 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_5 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_5 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_5 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_5 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_5 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_5 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_5 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_5 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_5 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_5 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_5 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_5 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_5 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_5 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_5 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_5 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_5 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_5 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_5 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_5 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_5 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_5 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_5 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_5 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_5 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_5 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_5 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_5 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_5 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_5 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_5 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_5 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_5 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_5 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_5 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_5 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_5 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_5 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_5 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_5 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_5 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_5 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_5 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_5 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_5 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_5 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_5 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_5 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_5 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_5 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_5 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_5 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_5 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_5 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_5 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_5 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_5 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_5 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_5 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_5 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_5 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_5 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_5 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_5 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_5 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_5 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_5 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_5 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_5 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_5 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_5 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_5 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_5 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_5 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_5 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_5 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_5 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_5 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_5 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_5 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_5 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_5 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_5 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_5 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_5 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_5 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_5 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_5 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_5 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_5 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_5 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_5 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_5 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_5 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_5 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_5 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_5 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_5 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_5 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_5 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_5 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_5 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_5 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_5 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_5 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_5 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_5 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_5 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_5 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_5 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_5 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_5 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_5 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_5 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_5 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_5 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_5 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_5 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_5 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_5 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_5 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_5 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_5 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_5 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_5 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_5 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_5 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_5 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_5 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_5 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_5 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_5 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_5 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_5 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_5 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_5 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_5 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_5 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_5 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_5 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_5 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_5 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_5 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_5 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_5 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_5 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_5 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_5 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_5 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_5 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_5 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_5 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_5 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_5 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_5 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_5 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_5 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_5 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_5 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_5 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_5 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_5 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_5 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_5 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_5 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_5 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_5 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_5 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_5 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_5 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_5 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_5 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_5 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_5 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_5 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_5 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_5 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_5 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_5 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_5 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_5 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_5 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_5 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_5 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_5 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_5 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_5 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_5 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_5 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_5 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_5 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_5 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_5 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_5 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_5 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_5 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_5 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_5 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_5 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_5 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_5 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_5 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_5 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_5 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_5 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_5 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_5 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_5 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_5 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_5 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_5 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_5 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_5 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_5 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_5 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_5 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_5 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_5 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_5 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_5 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_5 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_5 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_5 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_5 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_5 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_5 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_5 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_5 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_5 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_5 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_5 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_5 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_5 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_5 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_5 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_5 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_5 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_5 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_5 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_5 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_5 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_5 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_5 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_5 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_5 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_5 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_5 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_5 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_5 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_5 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_5 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_5 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_5 = sboxRom_254;
      default : _zz__zz_stateReg_5 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_9_1)
      8'b00000000 : _zz__zz_stateReg_9 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_9 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_9 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_9 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_9 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_9 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_9 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_9 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_9 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_9 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_9 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_9 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_9 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_9 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_9 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_9 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_9 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_9 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_9 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_9 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_9 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_9 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_9 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_9 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_9 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_9 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_9 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_9 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_9 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_9 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_9 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_9 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_9 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_9 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_9 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_9 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_9 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_9 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_9 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_9 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_9 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_9 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_9 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_9 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_9 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_9 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_9 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_9 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_9 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_9 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_9 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_9 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_9 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_9 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_9 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_9 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_9 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_9 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_9 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_9 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_9 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_9 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_9 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_9 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_9 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_9 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_9 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_9 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_9 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_9 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_9 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_9 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_9 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_9 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_9 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_9 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_9 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_9 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_9 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_9 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_9 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_9 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_9 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_9 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_9 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_9 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_9 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_9 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_9 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_9 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_9 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_9 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_9 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_9 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_9 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_9 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_9 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_9 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_9 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_9 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_9 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_9 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_9 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_9 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_9 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_9 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_9 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_9 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_9 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_9 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_9 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_9 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_9 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_9 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_9 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_9 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_9 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_9 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_9 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_9 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_9 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_9 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_9 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_9 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_9 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_9 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_9 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_9 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_9 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_9 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_9 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_9 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_9 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_9 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_9 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_9 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_9 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_9 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_9 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_9 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_9 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_9 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_9 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_9 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_9 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_9 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_9 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_9 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_9 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_9 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_9 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_9 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_9 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_9 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_9 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_9 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_9 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_9 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_9 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_9 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_9 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_9 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_9 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_9 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_9 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_9 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_9 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_9 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_9 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_9 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_9 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_9 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_9 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_9 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_9 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_9 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_9 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_9 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_9 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_9 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_9 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_9 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_9 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_9 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_9 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_9 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_9 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_9 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_9 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_9 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_9 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_9 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_9 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_9 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_9 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_9 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_9 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_9 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_9 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_9 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_9 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_9 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_9 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_9 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_9 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_9 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_9 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_9 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_9 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_9 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_9 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_9 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_9 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_9 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_9 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_9 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_9 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_9 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_9 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_9 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_9 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_9 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_9 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_9 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_9 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_9 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_9 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_9 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_9 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_9 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_9 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_9 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_9 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_9 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_9 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_9 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_9 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_9 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_9 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_9 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_9 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_9 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_9 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_9 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_9 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_9 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_9 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_9 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_9 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_9 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_9 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_9 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_9 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_9 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_9 = sboxRom_254;
      default : _zz__zz_stateReg_9 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_13_1)
      8'b00000000 : _zz__zz_stateReg_13 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_13 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_13 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_13 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_13 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_13 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_13 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_13 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_13 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_13 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_13 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_13 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_13 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_13 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_13 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_13 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_13 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_13 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_13 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_13 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_13 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_13 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_13 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_13 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_13 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_13 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_13 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_13 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_13 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_13 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_13 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_13 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_13 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_13 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_13 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_13 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_13 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_13 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_13 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_13 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_13 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_13 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_13 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_13 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_13 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_13 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_13 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_13 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_13 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_13 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_13 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_13 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_13 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_13 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_13 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_13 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_13 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_13 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_13 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_13 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_13 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_13 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_13 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_13 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_13 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_13 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_13 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_13 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_13 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_13 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_13 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_13 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_13 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_13 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_13 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_13 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_13 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_13 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_13 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_13 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_13 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_13 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_13 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_13 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_13 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_13 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_13 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_13 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_13 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_13 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_13 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_13 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_13 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_13 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_13 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_13 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_13 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_13 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_13 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_13 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_13 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_13 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_13 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_13 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_13 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_13 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_13 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_13 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_13 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_13 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_13 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_13 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_13 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_13 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_13 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_13 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_13 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_13 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_13 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_13 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_13 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_13 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_13 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_13 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_13 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_13 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_13 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_13 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_13 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_13 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_13 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_13 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_13 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_13 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_13 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_13 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_13 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_13 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_13 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_13 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_13 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_13 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_13 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_13 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_13 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_13 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_13 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_13 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_13 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_13 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_13 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_13 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_13 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_13 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_13 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_13 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_13 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_13 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_13 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_13 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_13 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_13 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_13 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_13 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_13 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_13 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_13 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_13 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_13 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_13 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_13 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_13 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_13 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_13 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_13 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_13 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_13 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_13 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_13 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_13 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_13 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_13 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_13 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_13 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_13 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_13 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_13 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_13 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_13 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_13 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_13 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_13 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_13 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_13 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_13 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_13 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_13 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_13 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_13 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_13 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_13 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_13 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_13 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_13 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_13 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_13 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_13 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_13 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_13 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_13 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_13 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_13 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_13 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_13 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_13 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_13 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_13 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_13 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_13 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_13 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_13 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_13 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_13 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_13 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_13 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_13 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_13 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_13 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_13 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_13 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_13 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_13 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_13 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_13 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_13 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_13 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_13 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_13 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_13 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_13 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_13 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_13 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_13 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_13 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_13 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_13 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_13 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_13 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_13 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_13 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_13 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_13 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_13 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_13 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_13 = sboxRom_254;
      default : _zz__zz_stateReg_13 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_17_1)
      8'b00000000 : _zz__zz_stateReg_17 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_17 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_17 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_17 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_17 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_17 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_17 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_17 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_17 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_17 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_17 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_17 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_17 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_17 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_17 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_17 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_17 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_17 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_17 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_17 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_17 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_17 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_17 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_17 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_17 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_17 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_17 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_17 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_17 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_17 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_17 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_17 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_17 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_17 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_17 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_17 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_17 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_17 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_17 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_17 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_17 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_17 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_17 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_17 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_17 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_17 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_17 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_17 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_17 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_17 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_17 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_17 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_17 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_17 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_17 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_17 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_17 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_17 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_17 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_17 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_17 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_17 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_17 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_17 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_17 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_17 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_17 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_17 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_17 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_17 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_17 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_17 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_17 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_17 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_17 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_17 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_17 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_17 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_17 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_17 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_17 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_17 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_17 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_17 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_17 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_17 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_17 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_17 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_17 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_17 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_17 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_17 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_17 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_17 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_17 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_17 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_17 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_17 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_17 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_17 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_17 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_17 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_17 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_17 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_17 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_17 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_17 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_17 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_17 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_17 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_17 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_17 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_17 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_17 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_17 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_17 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_17 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_17 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_17 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_17 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_17 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_17 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_17 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_17 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_17 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_17 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_17 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_17 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_17 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_17 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_17 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_17 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_17 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_17 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_17 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_17 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_17 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_17 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_17 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_17 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_17 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_17 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_17 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_17 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_17 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_17 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_17 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_17 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_17 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_17 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_17 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_17 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_17 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_17 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_17 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_17 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_17 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_17 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_17 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_17 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_17 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_17 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_17 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_17 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_17 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_17 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_17 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_17 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_17 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_17 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_17 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_17 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_17 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_17 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_17 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_17 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_17 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_17 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_17 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_17 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_17 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_17 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_17 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_17 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_17 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_17 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_17 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_17 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_17 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_17 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_17 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_17 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_17 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_17 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_17 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_17 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_17 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_17 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_17 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_17 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_17 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_17 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_17 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_17 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_17 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_17 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_17 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_17 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_17 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_17 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_17 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_17 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_17 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_17 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_17 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_17 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_17 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_17 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_17 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_17 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_17 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_17 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_17 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_17 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_17 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_17 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_17 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_17 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_17 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_17 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_17 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_17 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_17 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_17 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_17 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_17 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_17 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_17 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_17 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_17 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_17 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_17 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_17 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_17 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_17 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_17 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_17 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_17 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_17 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_17 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_17 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_17 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_17 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_17 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_17 = sboxRom_254;
      default : _zz__zz_stateReg_17 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_6_1)
      8'b00000000 : _zz__zz_stateReg_6 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_6 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_6 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_6 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_6 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_6 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_6 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_6 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_6 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_6 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_6 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_6 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_6 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_6 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_6 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_6 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_6 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_6 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_6 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_6 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_6 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_6 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_6 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_6 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_6 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_6 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_6 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_6 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_6 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_6 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_6 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_6 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_6 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_6 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_6 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_6 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_6 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_6 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_6 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_6 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_6 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_6 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_6 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_6 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_6 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_6 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_6 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_6 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_6 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_6 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_6 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_6 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_6 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_6 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_6 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_6 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_6 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_6 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_6 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_6 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_6 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_6 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_6 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_6 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_6 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_6 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_6 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_6 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_6 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_6 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_6 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_6 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_6 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_6 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_6 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_6 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_6 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_6 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_6 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_6 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_6 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_6 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_6 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_6 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_6 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_6 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_6 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_6 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_6 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_6 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_6 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_6 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_6 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_6 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_6 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_6 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_6 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_6 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_6 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_6 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_6 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_6 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_6 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_6 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_6 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_6 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_6 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_6 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_6 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_6 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_6 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_6 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_6 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_6 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_6 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_6 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_6 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_6 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_6 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_6 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_6 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_6 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_6 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_6 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_6 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_6 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_6 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_6 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_6 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_6 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_6 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_6 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_6 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_6 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_6 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_6 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_6 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_6 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_6 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_6 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_6 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_6 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_6 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_6 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_6 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_6 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_6 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_6 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_6 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_6 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_6 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_6 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_6 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_6 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_6 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_6 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_6 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_6 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_6 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_6 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_6 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_6 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_6 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_6 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_6 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_6 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_6 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_6 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_6 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_6 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_6 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_6 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_6 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_6 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_6 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_6 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_6 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_6 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_6 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_6 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_6 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_6 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_6 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_6 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_6 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_6 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_6 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_6 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_6 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_6 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_6 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_6 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_6 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_6 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_6 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_6 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_6 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_6 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_6 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_6 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_6 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_6 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_6 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_6 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_6 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_6 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_6 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_6 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_6 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_6 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_6 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_6 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_6 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_6 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_6 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_6 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_6 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_6 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_6 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_6 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_6 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_6 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_6 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_6 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_6 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_6 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_6 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_6 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_6 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_6 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_6 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_6 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_6 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_6 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_6 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_6 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_6 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_6 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_6 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_6 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_6 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_6 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_6 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_6 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_6 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_6 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_6 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_6 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_6 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_6 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_6 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_6 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_6 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_6 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_6 = sboxRom_254;
      default : _zz__zz_stateReg_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_10_1)
      8'b00000000 : _zz__zz_stateReg_10 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_10 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_10 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_10 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_10 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_10 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_10 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_10 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_10 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_10 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_10 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_10 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_10 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_10 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_10 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_10 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_10 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_10 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_10 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_10 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_10 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_10 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_10 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_10 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_10 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_10 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_10 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_10 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_10 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_10 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_10 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_10 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_10 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_10 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_10 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_10 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_10 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_10 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_10 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_10 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_10 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_10 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_10 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_10 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_10 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_10 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_10 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_10 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_10 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_10 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_10 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_10 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_10 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_10 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_10 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_10 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_10 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_10 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_10 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_10 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_10 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_10 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_10 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_10 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_10 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_10 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_10 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_10 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_10 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_10 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_10 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_10 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_10 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_10 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_10 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_10 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_10 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_10 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_10 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_10 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_10 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_10 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_10 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_10 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_10 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_10 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_10 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_10 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_10 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_10 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_10 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_10 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_10 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_10 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_10 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_10 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_10 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_10 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_10 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_10 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_10 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_10 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_10 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_10 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_10 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_10 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_10 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_10 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_10 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_10 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_10 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_10 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_10 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_10 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_10 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_10 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_10 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_10 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_10 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_10 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_10 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_10 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_10 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_10 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_10 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_10 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_10 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_10 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_10 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_10 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_10 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_10 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_10 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_10 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_10 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_10 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_10 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_10 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_10 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_10 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_10 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_10 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_10 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_10 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_10 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_10 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_10 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_10 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_10 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_10 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_10 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_10 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_10 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_10 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_10 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_10 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_10 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_10 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_10 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_10 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_10 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_10 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_10 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_10 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_10 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_10 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_10 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_10 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_10 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_10 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_10 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_10 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_10 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_10 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_10 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_10 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_10 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_10 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_10 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_10 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_10 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_10 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_10 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_10 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_10 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_10 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_10 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_10 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_10 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_10 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_10 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_10 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_10 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_10 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_10 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_10 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_10 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_10 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_10 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_10 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_10 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_10 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_10 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_10 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_10 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_10 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_10 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_10 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_10 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_10 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_10 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_10 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_10 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_10 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_10 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_10 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_10 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_10 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_10 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_10 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_10 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_10 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_10 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_10 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_10 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_10 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_10 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_10 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_10 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_10 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_10 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_10 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_10 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_10 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_10 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_10 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_10 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_10 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_10 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_10 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_10 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_10 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_10 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_10 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_10 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_10 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_10 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_10 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_10 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_10 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_10 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_10 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_10 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_10 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_10 = sboxRom_254;
      default : _zz__zz_stateReg_10 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_14_1)
      8'b00000000 : _zz__zz_stateReg_14 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_14 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_14 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_14 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_14 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_14 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_14 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_14 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_14 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_14 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_14 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_14 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_14 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_14 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_14 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_14 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_14 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_14 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_14 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_14 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_14 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_14 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_14 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_14 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_14 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_14 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_14 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_14 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_14 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_14 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_14 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_14 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_14 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_14 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_14 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_14 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_14 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_14 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_14 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_14 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_14 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_14 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_14 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_14 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_14 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_14 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_14 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_14 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_14 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_14 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_14 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_14 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_14 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_14 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_14 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_14 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_14 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_14 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_14 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_14 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_14 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_14 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_14 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_14 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_14 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_14 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_14 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_14 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_14 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_14 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_14 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_14 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_14 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_14 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_14 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_14 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_14 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_14 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_14 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_14 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_14 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_14 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_14 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_14 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_14 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_14 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_14 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_14 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_14 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_14 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_14 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_14 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_14 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_14 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_14 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_14 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_14 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_14 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_14 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_14 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_14 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_14 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_14 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_14 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_14 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_14 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_14 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_14 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_14 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_14 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_14 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_14 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_14 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_14 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_14 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_14 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_14 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_14 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_14 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_14 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_14 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_14 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_14 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_14 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_14 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_14 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_14 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_14 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_14 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_14 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_14 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_14 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_14 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_14 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_14 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_14 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_14 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_14 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_14 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_14 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_14 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_14 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_14 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_14 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_14 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_14 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_14 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_14 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_14 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_14 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_14 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_14 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_14 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_14 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_14 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_14 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_14 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_14 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_14 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_14 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_14 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_14 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_14 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_14 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_14 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_14 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_14 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_14 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_14 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_14 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_14 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_14 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_14 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_14 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_14 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_14 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_14 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_14 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_14 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_14 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_14 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_14 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_14 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_14 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_14 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_14 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_14 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_14 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_14 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_14 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_14 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_14 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_14 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_14 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_14 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_14 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_14 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_14 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_14 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_14 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_14 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_14 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_14 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_14 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_14 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_14 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_14 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_14 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_14 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_14 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_14 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_14 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_14 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_14 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_14 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_14 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_14 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_14 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_14 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_14 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_14 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_14 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_14 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_14 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_14 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_14 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_14 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_14 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_14 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_14 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_14 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_14 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_14 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_14 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_14 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_14 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_14 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_14 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_14 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_14 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_14 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_14 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_14 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_14 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_14 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_14 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_14 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_14 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_14 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_14 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_14 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_14 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_14 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_14 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_14 = sboxRom_254;
      default : _zz__zz_stateReg_14 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_18_1)
      8'b00000000 : _zz__zz_stateReg_18 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_18 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_18 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_18 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_18 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_18 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_18 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_18 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_18 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_18 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_18 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_18 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_18 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_18 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_18 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_18 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_18 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_18 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_18 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_18 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_18 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_18 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_18 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_18 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_18 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_18 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_18 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_18 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_18 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_18 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_18 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_18 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_18 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_18 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_18 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_18 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_18 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_18 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_18 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_18 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_18 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_18 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_18 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_18 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_18 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_18 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_18 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_18 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_18 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_18 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_18 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_18 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_18 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_18 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_18 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_18 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_18 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_18 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_18 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_18 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_18 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_18 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_18 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_18 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_18 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_18 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_18 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_18 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_18 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_18 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_18 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_18 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_18 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_18 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_18 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_18 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_18 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_18 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_18 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_18 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_18 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_18 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_18 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_18 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_18 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_18 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_18 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_18 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_18 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_18 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_18 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_18 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_18 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_18 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_18 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_18 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_18 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_18 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_18 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_18 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_18 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_18 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_18 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_18 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_18 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_18 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_18 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_18 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_18 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_18 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_18 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_18 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_18 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_18 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_18 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_18 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_18 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_18 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_18 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_18 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_18 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_18 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_18 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_18 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_18 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_18 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_18 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_18 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_18 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_18 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_18 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_18 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_18 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_18 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_18 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_18 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_18 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_18 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_18 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_18 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_18 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_18 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_18 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_18 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_18 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_18 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_18 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_18 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_18 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_18 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_18 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_18 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_18 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_18 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_18 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_18 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_18 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_18 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_18 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_18 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_18 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_18 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_18 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_18 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_18 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_18 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_18 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_18 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_18 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_18 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_18 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_18 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_18 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_18 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_18 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_18 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_18 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_18 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_18 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_18 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_18 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_18 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_18 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_18 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_18 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_18 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_18 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_18 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_18 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_18 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_18 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_18 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_18 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_18 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_18 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_18 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_18 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_18 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_18 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_18 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_18 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_18 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_18 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_18 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_18 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_18 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_18 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_18 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_18 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_18 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_18 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_18 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_18 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_18 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_18 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_18 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_18 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_18 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_18 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_18 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_18 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_18 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_18 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_18 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_18 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_18 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_18 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_18 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_18 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_18 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_18 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_18 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_18 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_18 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_18 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_18 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_18 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_18 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_18 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_18 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_18 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_18 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_18 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_18 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_18 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_18 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_18 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_18 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_18 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_18 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_18 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_18 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_18 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_18 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_18 = sboxRom_254;
      default : _zz__zz_stateReg_18 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_7_1)
      8'b00000000 : _zz__zz_stateReg_7 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_7 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_7 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_7 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_7 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_7 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_7 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_7 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_7 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_7 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_7 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_7 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_7 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_7 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_7 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_7 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_7 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_7 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_7 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_7 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_7 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_7 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_7 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_7 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_7 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_7 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_7 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_7 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_7 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_7 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_7 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_7 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_7 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_7 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_7 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_7 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_7 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_7 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_7 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_7 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_7 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_7 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_7 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_7 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_7 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_7 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_7 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_7 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_7 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_7 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_7 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_7 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_7 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_7 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_7 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_7 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_7 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_7 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_7 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_7 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_7 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_7 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_7 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_7 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_7 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_7 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_7 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_7 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_7 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_7 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_7 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_7 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_7 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_7 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_7 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_7 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_7 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_7 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_7 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_7 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_7 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_7 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_7 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_7 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_7 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_7 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_7 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_7 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_7 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_7 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_7 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_7 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_7 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_7 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_7 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_7 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_7 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_7 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_7 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_7 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_7 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_7 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_7 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_7 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_7 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_7 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_7 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_7 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_7 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_7 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_7 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_7 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_7 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_7 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_7 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_7 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_7 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_7 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_7 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_7 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_7 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_7 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_7 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_7 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_7 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_7 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_7 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_7 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_7 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_7 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_7 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_7 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_7 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_7 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_7 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_7 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_7 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_7 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_7 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_7 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_7 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_7 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_7 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_7 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_7 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_7 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_7 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_7 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_7 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_7 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_7 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_7 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_7 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_7 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_7 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_7 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_7 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_7 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_7 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_7 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_7 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_7 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_7 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_7 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_7 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_7 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_7 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_7 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_7 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_7 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_7 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_7 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_7 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_7 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_7 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_7 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_7 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_7 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_7 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_7 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_7 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_7 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_7 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_7 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_7 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_7 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_7 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_7 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_7 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_7 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_7 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_7 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_7 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_7 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_7 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_7 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_7 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_7 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_7 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_7 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_7 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_7 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_7 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_7 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_7 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_7 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_7 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_7 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_7 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_7 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_7 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_7 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_7 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_7 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_7 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_7 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_7 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_7 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_7 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_7 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_7 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_7 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_7 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_7 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_7 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_7 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_7 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_7 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_7 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_7 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_7 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_7 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_7 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_7 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_7 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_7 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_7 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_7 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_7 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_7 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_7 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_7 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_7 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_7 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_7 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_7 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_7 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_7 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_7 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_7 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_7 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_7 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_7 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_7 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_7 = sboxRom_254;
      default : _zz__zz_stateReg_7 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_11_1)
      8'b00000000 : _zz__zz_stateReg_11 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_11 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_11 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_11 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_11 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_11 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_11 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_11 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_11 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_11 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_11 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_11 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_11 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_11 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_11 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_11 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_11 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_11 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_11 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_11 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_11 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_11 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_11 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_11 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_11 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_11 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_11 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_11 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_11 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_11 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_11 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_11 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_11 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_11 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_11 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_11 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_11 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_11 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_11 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_11 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_11 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_11 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_11 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_11 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_11 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_11 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_11 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_11 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_11 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_11 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_11 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_11 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_11 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_11 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_11 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_11 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_11 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_11 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_11 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_11 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_11 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_11 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_11 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_11 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_11 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_11 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_11 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_11 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_11 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_11 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_11 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_11 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_11 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_11 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_11 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_11 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_11 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_11 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_11 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_11 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_11 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_11 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_11 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_11 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_11 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_11 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_11 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_11 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_11 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_11 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_11 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_11 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_11 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_11 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_11 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_11 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_11 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_11 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_11 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_11 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_11 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_11 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_11 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_11 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_11 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_11 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_11 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_11 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_11 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_11 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_11 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_11 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_11 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_11 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_11 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_11 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_11 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_11 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_11 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_11 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_11 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_11 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_11 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_11 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_11 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_11 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_11 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_11 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_11 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_11 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_11 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_11 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_11 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_11 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_11 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_11 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_11 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_11 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_11 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_11 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_11 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_11 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_11 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_11 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_11 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_11 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_11 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_11 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_11 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_11 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_11 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_11 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_11 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_11 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_11 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_11 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_11 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_11 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_11 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_11 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_11 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_11 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_11 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_11 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_11 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_11 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_11 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_11 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_11 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_11 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_11 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_11 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_11 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_11 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_11 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_11 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_11 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_11 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_11 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_11 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_11 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_11 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_11 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_11 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_11 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_11 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_11 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_11 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_11 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_11 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_11 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_11 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_11 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_11 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_11 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_11 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_11 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_11 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_11 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_11 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_11 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_11 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_11 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_11 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_11 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_11 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_11 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_11 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_11 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_11 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_11 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_11 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_11 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_11 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_11 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_11 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_11 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_11 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_11 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_11 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_11 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_11 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_11 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_11 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_11 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_11 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_11 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_11 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_11 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_11 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_11 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_11 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_11 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_11 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_11 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_11 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_11 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_11 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_11 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_11 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_11 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_11 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_11 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_11 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_11 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_11 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_11 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_11 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_11 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_11 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_11 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_11 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_11 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_11 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_11 = sboxRom_254;
      default : _zz__zz_stateReg_11 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_15_1)
      8'b00000000 : _zz__zz_stateReg_15 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_15 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_15 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_15 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_15 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_15 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_15 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_15 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_15 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_15 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_15 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_15 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_15 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_15 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_15 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_15 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_15 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_15 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_15 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_15 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_15 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_15 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_15 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_15 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_15 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_15 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_15 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_15 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_15 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_15 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_15 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_15 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_15 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_15 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_15 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_15 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_15 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_15 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_15 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_15 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_15 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_15 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_15 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_15 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_15 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_15 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_15 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_15 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_15 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_15 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_15 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_15 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_15 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_15 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_15 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_15 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_15 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_15 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_15 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_15 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_15 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_15 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_15 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_15 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_15 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_15 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_15 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_15 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_15 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_15 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_15 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_15 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_15 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_15 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_15 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_15 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_15 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_15 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_15 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_15 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_15 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_15 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_15 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_15 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_15 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_15 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_15 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_15 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_15 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_15 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_15 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_15 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_15 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_15 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_15 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_15 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_15 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_15 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_15 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_15 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_15 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_15 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_15 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_15 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_15 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_15 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_15 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_15 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_15 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_15 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_15 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_15 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_15 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_15 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_15 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_15 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_15 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_15 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_15 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_15 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_15 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_15 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_15 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_15 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_15 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_15 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_15 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_15 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_15 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_15 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_15 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_15 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_15 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_15 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_15 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_15 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_15 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_15 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_15 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_15 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_15 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_15 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_15 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_15 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_15 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_15 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_15 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_15 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_15 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_15 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_15 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_15 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_15 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_15 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_15 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_15 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_15 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_15 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_15 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_15 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_15 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_15 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_15 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_15 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_15 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_15 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_15 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_15 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_15 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_15 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_15 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_15 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_15 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_15 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_15 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_15 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_15 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_15 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_15 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_15 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_15 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_15 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_15 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_15 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_15 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_15 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_15 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_15 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_15 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_15 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_15 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_15 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_15 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_15 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_15 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_15 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_15 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_15 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_15 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_15 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_15 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_15 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_15 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_15 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_15 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_15 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_15 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_15 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_15 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_15 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_15 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_15 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_15 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_15 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_15 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_15 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_15 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_15 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_15 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_15 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_15 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_15 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_15 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_15 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_15 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_15 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_15 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_15 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_15 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_15 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_15 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_15 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_15 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_15 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_15 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_15 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_15 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_15 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_15 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_15 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_15 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_15 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_15 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_15 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_15 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_15 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_15 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_15 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_15 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_15 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_15 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_15 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_15 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_15 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_15 = sboxRom_254;
      default : _zz__zz_stateReg_15 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_19_1)
      8'b00000000 : _zz__zz_stateReg_19 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_19 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_19 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_19 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_19 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_19 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_19 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_19 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_19 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_19 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_19 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_19 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_19 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_19 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_19 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_19 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_19 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_19 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_19 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_19 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_19 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_19 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_19 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_19 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_19 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_19 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_19 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_19 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_19 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_19 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_19 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_19 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_19 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_19 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_19 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_19 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_19 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_19 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_19 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_19 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_19 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_19 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_19 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_19 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_19 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_19 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_19 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_19 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_19 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_19 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_19 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_19 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_19 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_19 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_19 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_19 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_19 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_19 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_19 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_19 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_19 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_19 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_19 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_19 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_19 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_19 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_19 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_19 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_19 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_19 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_19 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_19 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_19 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_19 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_19 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_19 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_19 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_19 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_19 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_19 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_19 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_19 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_19 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_19 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_19 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_19 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_19 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_19 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_19 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_19 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_19 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_19 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_19 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_19 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_19 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_19 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_19 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_19 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_19 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_19 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_19 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_19 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_19 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_19 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_19 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_19 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_19 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_19 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_19 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_19 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_19 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_19 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_19 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_19 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_19 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_19 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_19 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_19 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_19 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_19 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_19 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_19 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_19 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_19 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_19 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_19 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_19 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_19 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_19 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_19 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_19 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_19 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_19 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_19 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_19 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_19 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_19 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_19 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_19 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_19 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_19 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_19 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_19 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_19 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_19 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_19 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_19 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_19 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_19 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_19 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_19 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_19 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_19 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_19 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_19 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_19 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_19 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_19 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_19 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_19 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_19 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_19 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_19 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_19 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_19 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_19 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_19 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_19 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_19 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_19 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_19 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_19 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_19 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_19 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_19 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_19 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_19 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_19 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_19 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_19 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_19 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_19 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_19 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_19 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_19 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_19 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_19 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_19 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_19 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_19 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_19 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_19 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_19 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_19 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_19 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_19 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_19 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_19 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_19 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_19 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_19 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_19 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_19 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_19 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_19 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_19 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_19 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_19 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_19 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_19 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_19 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_19 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_19 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_19 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_19 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_19 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_19 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_19 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_19 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_19 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_19 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_19 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_19 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_19 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_19 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_19 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_19 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_19 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_19 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_19 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_19 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_19 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_19 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_19 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_19 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_19 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_19 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_19 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_19 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_19 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_19 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_19 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_19 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_19 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_19 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_19 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_19 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_19 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_19 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_19 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_19 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_19 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_19 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_19 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_19 = sboxRom_254;
      default : _zz__zz_stateReg_19 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(rconCounter)
      4'b0000 : _zz__zz_roundKeyReg_0 = rcon_0;
      4'b0001 : _zz__zz_roundKeyReg_0 = rcon_1;
      4'b0010 : _zz__zz_roundKeyReg_0 = rcon_2;
      4'b0011 : _zz__zz_roundKeyReg_0 = rcon_3;
      4'b0100 : _zz__zz_roundKeyReg_0 = rcon_4;
      4'b0101 : _zz__zz_roundKeyReg_0 = rcon_5;
      4'b0110 : _zz__zz_roundKeyReg_0 = rcon_6;
      4'b0111 : _zz__zz_roundKeyReg_0 = rcon_7;
      4'b1000 : _zz__zz_roundKeyReg_0 = rcon_8;
      default : _zz__zz_roundKeyReg_0 = rcon_9;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_1)
      8'b00000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_3)
      8'b00000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_5)
      8'b00000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2_4 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_2_7)
      8'b00000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_2_6 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_2_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_1)
      8'b00000000 : _zz__zz_stateReg_71 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71 = sboxRom_254;
      default : _zz__zz_stateReg_71 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_3)
      8'b00000000 : _zz__zz_stateReg_71_2 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71_2 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71_2 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71_2 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71_2 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71_2 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71_2 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71_2 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71_2 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71_2 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71_2 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71_2 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71_2 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71_2 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71_2 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71_2 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71_2 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71_2 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71_2 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71_2 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71_2 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71_2 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71_2 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71_2 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71_2 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71_2 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71_2 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71_2 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71_2 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71_2 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71_2 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71_2 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71_2 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71_2 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71_2 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71_2 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71_2 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71_2 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71_2 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71_2 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71_2 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71_2 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71_2 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71_2 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71_2 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71_2 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71_2 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71_2 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71_2 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71_2 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71_2 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71_2 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71_2 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71_2 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71_2 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71_2 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71_2 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71_2 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71_2 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71_2 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71_2 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71_2 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71_2 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71_2 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71_2 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71_2 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71_2 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71_2 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71_2 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71_2 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71_2 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71_2 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71_2 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71_2 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71_2 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71_2 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71_2 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71_2 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71_2 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71_2 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71_2 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71_2 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71_2 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71_2 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71_2 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71_2 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71_2 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71_2 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71_2 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71_2 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71_2 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71_2 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71_2 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71_2 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71_2 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71_2 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71_2 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71_2 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71_2 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71_2 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71_2 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71_2 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71_2 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71_2 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71_2 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71_2 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71_2 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71_2 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71_2 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71_2 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71_2 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71_2 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71_2 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71_2 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71_2 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71_2 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71_2 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71_2 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71_2 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71_2 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71_2 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71_2 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71_2 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71_2 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71_2 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71_2 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71_2 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71_2 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71_2 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71_2 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71_2 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71_2 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71_2 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71_2 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71_2 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71_2 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71_2 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71_2 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71_2 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71_2 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71_2 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71_2 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71_2 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71_2 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71_2 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71_2 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71_2 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71_2 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71_2 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71_2 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71_2 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71_2 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71_2 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71_2 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71_2 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71_2 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71_2 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71_2 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71_2 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71_2 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71_2 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71_2 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71_2 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71_2 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71_2 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71_2 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71_2 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71_2 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71_2 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71_2 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71_2 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71_2 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71_2 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71_2 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71_2 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71_2 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71_2 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71_2 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71_2 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71_2 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71_2 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71_2 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71_2 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71_2 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71_2 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71_2 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71_2 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71_2 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71_2 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71_2 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71_2 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71_2 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71_2 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71_2 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71_2 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71_2 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71_2 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71_2 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71_2 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71_2 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71_2 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71_2 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71_2 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71_2 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71_2 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71_2 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71_2 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71_2 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71_2 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71_2 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71_2 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71_2 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71_2 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71_2 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71_2 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71_2 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71_2 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71_2 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71_2 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71_2 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71_2 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71_2 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71_2 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71_2 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71_2 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71_2 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71_2 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71_2 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71_2 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71_2 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71_2 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71_2 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71_2 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71_2 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71_2 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71_2 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71_2 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71_2 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71_2 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71_2 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71_2 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71_2 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71_2 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71_2 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71_2 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71_2 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71_2 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71_2 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71_2 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71_2 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71_2 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71_2 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71_2 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71_2 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71_2 = sboxRom_254;
      default : _zz__zz_stateReg_71_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_5)
      8'b00000000 : _zz__zz_stateReg_71_4 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71_4 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71_4 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71_4 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71_4 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71_4 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71_4 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71_4 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71_4 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71_4 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71_4 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71_4 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71_4 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71_4 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71_4 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71_4 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71_4 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71_4 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71_4 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71_4 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71_4 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71_4 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71_4 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71_4 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71_4 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71_4 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71_4 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71_4 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71_4 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71_4 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71_4 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71_4 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71_4 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71_4 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71_4 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71_4 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71_4 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71_4 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71_4 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71_4 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71_4 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71_4 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71_4 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71_4 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71_4 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71_4 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71_4 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71_4 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71_4 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71_4 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71_4 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71_4 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71_4 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71_4 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71_4 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71_4 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71_4 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71_4 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71_4 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71_4 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71_4 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71_4 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71_4 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71_4 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71_4 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71_4 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71_4 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71_4 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71_4 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71_4 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71_4 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71_4 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71_4 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71_4 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71_4 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71_4 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71_4 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71_4 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71_4 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71_4 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71_4 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71_4 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71_4 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71_4 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71_4 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71_4 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71_4 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71_4 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71_4 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71_4 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71_4 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71_4 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71_4 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71_4 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71_4 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71_4 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71_4 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71_4 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71_4 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71_4 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71_4 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71_4 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71_4 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71_4 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71_4 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71_4 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71_4 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71_4 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71_4 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71_4 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71_4 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71_4 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71_4 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71_4 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71_4 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71_4 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71_4 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71_4 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71_4 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71_4 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71_4 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71_4 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71_4 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71_4 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71_4 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71_4 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71_4 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71_4 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71_4 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71_4 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71_4 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71_4 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71_4 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71_4 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71_4 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71_4 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71_4 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71_4 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71_4 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71_4 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71_4 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71_4 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71_4 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71_4 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71_4 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71_4 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71_4 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71_4 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71_4 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71_4 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71_4 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71_4 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71_4 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71_4 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71_4 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71_4 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71_4 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71_4 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71_4 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71_4 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71_4 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71_4 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71_4 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71_4 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71_4 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71_4 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71_4 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71_4 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71_4 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71_4 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71_4 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71_4 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71_4 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71_4 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71_4 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71_4 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71_4 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71_4 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71_4 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71_4 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71_4 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71_4 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71_4 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71_4 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71_4 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71_4 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71_4 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71_4 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71_4 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71_4 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71_4 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71_4 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71_4 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71_4 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71_4 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71_4 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71_4 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71_4 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71_4 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71_4 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71_4 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71_4 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71_4 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71_4 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71_4 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71_4 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71_4 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71_4 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71_4 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71_4 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71_4 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71_4 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71_4 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71_4 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71_4 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71_4 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71_4 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71_4 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71_4 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71_4 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71_4 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71_4 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71_4 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71_4 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71_4 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71_4 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71_4 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71_4 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71_4 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71_4 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71_4 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71_4 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71_4 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71_4 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71_4 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71_4 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71_4 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71_4 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71_4 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71_4 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71_4 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71_4 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71_4 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71_4 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71_4 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71_4 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71_4 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71_4 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71_4 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71_4 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71_4 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71_4 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71_4 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71_4 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71_4 = sboxRom_254;
      default : _zz__zz_stateReg_71_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_71_7)
      8'b00000000 : _zz__zz_stateReg_71_6 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_71_6 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_71_6 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_71_6 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_71_6 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_71_6 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_71_6 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_71_6 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_71_6 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_71_6 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_71_6 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_71_6 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_71_6 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_71_6 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_71_6 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_71_6 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_71_6 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_71_6 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_71_6 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_71_6 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_71_6 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_71_6 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_71_6 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_71_6 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_71_6 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_71_6 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_71_6 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_71_6 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_71_6 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_71_6 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_71_6 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_71_6 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_71_6 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_71_6 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_71_6 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_71_6 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_71_6 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_71_6 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_71_6 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_71_6 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_71_6 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_71_6 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_71_6 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_71_6 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_71_6 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_71_6 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_71_6 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_71_6 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_71_6 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_71_6 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_71_6 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_71_6 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_71_6 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_71_6 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_71_6 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_71_6 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_71_6 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_71_6 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_71_6 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_71_6 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_71_6 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_71_6 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_71_6 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_71_6 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_71_6 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_71_6 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_71_6 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_71_6 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_71_6 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_71_6 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_71_6 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_71_6 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_71_6 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_71_6 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_71_6 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_71_6 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_71_6 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_71_6 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_71_6 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_71_6 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_71_6 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_71_6 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_71_6 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_71_6 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_71_6 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_71_6 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_71_6 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_71_6 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_71_6 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_71_6 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_71_6 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_71_6 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_71_6 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_71_6 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_71_6 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_71_6 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_71_6 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_71_6 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_71_6 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_71_6 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_71_6 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_71_6 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_71_6 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_71_6 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_71_6 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_71_6 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_71_6 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_71_6 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_71_6 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_71_6 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_71_6 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_71_6 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_71_6 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_71_6 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_71_6 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_71_6 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_71_6 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_71_6 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_71_6 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_71_6 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_71_6 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_71_6 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_71_6 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_71_6 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_71_6 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_71_6 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_71_6 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_71_6 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_71_6 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_71_6 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_71_6 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_71_6 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_71_6 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_71_6 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_71_6 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_71_6 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_71_6 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_71_6 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_71_6 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_71_6 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_71_6 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_71_6 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_71_6 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_71_6 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_71_6 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_71_6 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_71_6 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_71_6 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_71_6 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_71_6 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_71_6 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_71_6 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_71_6 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_71_6 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_71_6 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_71_6 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_71_6 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_71_6 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_71_6 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_71_6 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_71_6 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_71_6 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_71_6 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_71_6 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_71_6 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_71_6 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_71_6 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_71_6 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_71_6 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_71_6 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_71_6 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_71_6 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_71_6 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_71_6 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_71_6 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_71_6 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_71_6 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_71_6 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_71_6 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_71_6 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_71_6 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_71_6 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_71_6 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_71_6 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_71_6 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_71_6 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_71_6 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_71_6 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_71_6 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_71_6 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_71_6 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_71_6 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_71_6 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_71_6 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_71_6 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_71_6 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_71_6 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_71_6 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_71_6 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_71_6 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_71_6 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_71_6 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_71_6 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_71_6 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_71_6 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_71_6 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_71_6 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_71_6 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_71_6 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_71_6 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_71_6 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_71_6 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_71_6 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_71_6 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_71_6 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_71_6 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_71_6 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_71_6 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_71_6 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_71_6 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_71_6 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_71_6 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_71_6 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_71_6 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_71_6 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_71_6 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_71_6 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_71_6 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_71_6 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_71_6 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_71_6 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_71_6 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_71_6 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_71_6 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_71_6 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_71_6 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_71_6 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_71_6 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_71_6 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_71_6 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_71_6 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_71_6 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_71_6 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_71_6 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_71_6 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_71_6 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_71_6 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_71_6 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_71_6 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_71_6 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_71_6 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_71_6 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_71_6 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_71_6 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_71_6 = sboxRom_254;
      default : _zz__zz_stateReg_71_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(precomputeCounter)
      4'b0000 : _zz__zz_stateReg_71_8 = rcon_0;
      4'b0001 : _zz__zz_stateReg_71_8 = rcon_1;
      4'b0010 : _zz__zz_stateReg_71_8 = rcon_2;
      4'b0011 : _zz__zz_stateReg_71_8 = rcon_3;
      4'b0100 : _zz__zz_stateReg_71_8 = rcon_4;
      4'b0101 : _zz__zz_stateReg_71_8 = rcon_5;
      4'b0110 : _zz__zz_stateReg_71_8 = rcon_6;
      4'b0111 : _zz__zz_stateReg_71_8 = rcon_7;
      4'b1000 : _zz__zz_stateReg_71_8 = rcon_8;
      default : _zz__zz_stateReg_71_8 = rcon_9;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_4_1)
      8'b00000000 : _zz__zz_roundKeyReg_0_4 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_4 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_4 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_4 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_4 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_4 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_4 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_4 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_4 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_4 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_4 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_4 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_4 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_4 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_4 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_4 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_4 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_4 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_4 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_4 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_4 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_4 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_4 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_4 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_4 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_4 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_4 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_4 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_4 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_4 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_4 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_4 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_4 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_4 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_4 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_4 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_4 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_4 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_4 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_4 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_4 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_4 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_4 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_4 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_4 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_4 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_4 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_4 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_4 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_4 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_4 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_4 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_4 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_4 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_4 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_4 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_4 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_4 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_4 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_4 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_4 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_4 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_4 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_4 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_4 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_4 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_4 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_4 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_4 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_4 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_4 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_4 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_4 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_4 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_4 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_4 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_4 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_4 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_4 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_4 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_4 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_4 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_4 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_4 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_4 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_4 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_4 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_4 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_4 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_4 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_4 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_4 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_4 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_4 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_4 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_4 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_4 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_4 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_4 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_4 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_4 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_4 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_4 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_4 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_4 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_4 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_4 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_4 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_4 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_4 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_4 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_4 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_4 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_4 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_4 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_4 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_4 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_4 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_4 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_4 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_4 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_4 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_4 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_4 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_4 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_4 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_4 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_4 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_4 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_4 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_4 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_4 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_4 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_4 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_4 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_4 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_4 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_4 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_4 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_4 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_4 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_4 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_4 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_4 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_4 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_4 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_4 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_4 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_4 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_4 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_4 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_4 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_4 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_4 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_4 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_4 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_4 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_4 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_4 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_4 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_4 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_4 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_4 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_4 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_4 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_4 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_4 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_4 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_4 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_4 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_4 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_4 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_4 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_4 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_4 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_4 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_4 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_4 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_4 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_4 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_4 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_4 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_4 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_4 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_4 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_4 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_4 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_4 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_4 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_4 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_4 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_4 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_4 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_4 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_4 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_4 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_4 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_4 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_4 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_4 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_4 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_4 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_4 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_4 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_4 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_4 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_4 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_4 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_4 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_4 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_4 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_4 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_4 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_4 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_4 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_4 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_4 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_4 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_4 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_4 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_4 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_4 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_4 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_4 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_4 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_4 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_4 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_4 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_4 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_4 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_4 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_4 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_4 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_4 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_4 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_4 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_4 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_4 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_4 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_4 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_4 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_4 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_4 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_4 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_4 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_4 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_4 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_4 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_4 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_4 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_4 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_4 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_4 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_4 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_4 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_4_3)
      8'b00000000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_4_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_4_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_4_5)
      8'b00000000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_4_4 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_4_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_4_7)
      8'b00000000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_4_6 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_4_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_3)
      8'b00000000 : _zz__zz_stateReg_75_2 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_2 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_2 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_2 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_2 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_2 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_2 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_2 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_2 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_2 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_2 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_2 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_2 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_2 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_2 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_2 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_2 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_2 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_2 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_2 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_2 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_2 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_2 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_2 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_2 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_2 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_2 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_2 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_2 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_2 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_2 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_2 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_2 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_2 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_2 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_2 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_2 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_2 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_2 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_2 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_2 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_2 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_2 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_2 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_2 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_2 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_2 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_2 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_2 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_2 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_2 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_2 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_2 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_2 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_2 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_2 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_2 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_2 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_2 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_2 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_2 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_2 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_2 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_2 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_2 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_2 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_2 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_2 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_2 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_2 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_2 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_2 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_2 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_2 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_2 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_2 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_2 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_2 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_2 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_2 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_2 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_2 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_2 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_2 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_2 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_2 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_2 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_2 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_2 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_2 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_2 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_2 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_2 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_2 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_2 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_2 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_2 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_2 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_2 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_2 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_2 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_2 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_2 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_2 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_2 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_2 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_2 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_2 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_2 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_2 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_2 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_2 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_2 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_2 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_2 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_2 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_2 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_2 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_2 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_2 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_2 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_2 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_2 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_2 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_2 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_2 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_2 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_2 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_2 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_2 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_2 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_2 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_2 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_2 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_2 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_2 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_2 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_2 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_2 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_2 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_2 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_2 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_2 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_2 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_2 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_2 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_2 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_2 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_2 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_2 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_2 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_2 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_2 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_2 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_2 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_2 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_2 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_2 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_2 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_2 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_2 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_2 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_2 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_2 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_2 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_2 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_2 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_2 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_2 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_2 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_2 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_2 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_2 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_2 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_2 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_2 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_2 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_2 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_2 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_2 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_2 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_2 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_2 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_2 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_2 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_2 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_2 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_2 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_2 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_2 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_2 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_2 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_2 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_2 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_2 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_2 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_2 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_2 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_2 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_2 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_2 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_2 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_2 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_2 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_2 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_2 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_2 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_2 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_2 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_2 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_2 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_2 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_2 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_2 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_2 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_2 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_2 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_2 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_2 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_2 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_2 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_2 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_2 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_2 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_2 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_2 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_2 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_2 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_2 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_2 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_2 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_2 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_2 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_2 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_2 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_2 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_2 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_2 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_2 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_2 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_2 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_2 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_2 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_2 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_2 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_2 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_2 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_2 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_2 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_2 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_2 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_2 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_2 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_2 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_2 = invSboxRom_254;
      default : _zz__zz_stateReg_75_2 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_5)
      8'b00000000 : _zz__zz_stateReg_75_4 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_4 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_4 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_4 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_4 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_4 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_4 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_4 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_4 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_4 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_4 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_4 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_4 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_4 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_4 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_4 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_4 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_4 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_4 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_4 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_4 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_4 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_4 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_4 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_4 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_4 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_4 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_4 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_4 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_4 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_4 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_4 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_4 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_4 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_4 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_4 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_4 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_4 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_4 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_4 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_4 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_4 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_4 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_4 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_4 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_4 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_4 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_4 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_4 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_4 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_4 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_4 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_4 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_4 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_4 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_4 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_4 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_4 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_4 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_4 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_4 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_4 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_4 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_4 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_4 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_4 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_4 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_4 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_4 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_4 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_4 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_4 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_4 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_4 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_4 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_4 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_4 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_4 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_4 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_4 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_4 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_4 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_4 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_4 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_4 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_4 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_4 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_4 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_4 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_4 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_4 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_4 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_4 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_4 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_4 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_4 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_4 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_4 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_4 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_4 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_4 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_4 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_4 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_4 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_4 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_4 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_4 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_4 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_4 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_4 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_4 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_4 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_4 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_4 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_4 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_4 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_4 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_4 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_4 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_4 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_4 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_4 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_4 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_4 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_4 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_4 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_4 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_4 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_4 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_4 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_4 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_4 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_4 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_4 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_4 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_4 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_4 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_4 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_4 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_4 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_4 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_4 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_4 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_4 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_4 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_4 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_4 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_4 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_4 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_4 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_4 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_4 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_4 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_4 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_4 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_4 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_4 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_4 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_4 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_4 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_4 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_4 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_4 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_4 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_4 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_4 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_4 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_4 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_4 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_4 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_4 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_4 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_4 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_4 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_4 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_4 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_4 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_4 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_4 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_4 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_4 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_4 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_4 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_4 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_4 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_4 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_4 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_4 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_4 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_4 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_4 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_4 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_4 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_4 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_4 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_4 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_4 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_4 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_4 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_4 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_4 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_4 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_4 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_4 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_4 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_4 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_4 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_4 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_4 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_4 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_4 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_4 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_4 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_4 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_4 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_4 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_4 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_4 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_4 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_4 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_4 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_4 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_4 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_4 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_4 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_4 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_4 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_4 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_4 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_4 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_4 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_4 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_4 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_4 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_4 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_4 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_4 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_4 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_4 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_4 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_4 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_4 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_4 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_4 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_4 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_4 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_4 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_4 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_4 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_4 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_4 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_4 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_4 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_4 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_4 = invSboxRom_254;
      default : _zz__zz_stateReg_75_4 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_7)
      8'b00000000 : _zz__zz_stateReg_75_6 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_6 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_6 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_6 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_6 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_6 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_6 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_6 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_6 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_6 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_6 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_6 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_6 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_6 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_6 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_6 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_6 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_6 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_6 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_6 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_6 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_6 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_6 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_6 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_6 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_6 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_6 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_6 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_6 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_6 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_6 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_6 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_6 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_6 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_6 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_6 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_6 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_6 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_6 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_6 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_6 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_6 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_6 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_6 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_6 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_6 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_6 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_6 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_6 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_6 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_6 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_6 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_6 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_6 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_6 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_6 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_6 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_6 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_6 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_6 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_6 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_6 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_6 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_6 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_6 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_6 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_6 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_6 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_6 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_6 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_6 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_6 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_6 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_6 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_6 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_6 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_6 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_6 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_6 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_6 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_6 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_6 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_6 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_6 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_6 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_6 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_6 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_6 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_6 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_6 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_6 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_6 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_6 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_6 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_6 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_6 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_6 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_6 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_6 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_6 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_6 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_6 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_6 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_6 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_6 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_6 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_6 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_6 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_6 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_6 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_6 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_6 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_6 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_6 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_6 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_6 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_6 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_6 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_6 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_6 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_6 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_6 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_6 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_6 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_6 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_6 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_6 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_6 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_6 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_6 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_6 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_6 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_6 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_6 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_6 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_6 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_6 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_6 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_6 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_6 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_6 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_6 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_6 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_6 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_6 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_6 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_6 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_6 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_6 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_6 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_6 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_6 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_6 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_6 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_6 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_6 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_6 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_6 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_6 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_6 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_6 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_6 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_6 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_6 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_6 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_6 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_6 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_6 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_6 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_6 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_6 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_6 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_6 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_6 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_6 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_6 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_6 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_6 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_6 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_6 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_6 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_6 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_6 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_6 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_6 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_6 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_6 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_6 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_6 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_6 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_6 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_6 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_6 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_6 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_6 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_6 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_6 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_6 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_6 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_6 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_6 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_6 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_6 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_6 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_6 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_6 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_6 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_6 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_6 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_6 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_6 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_6 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_6 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_6 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_6 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_6 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_6 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_6 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_6 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_6 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_6 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_6 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_6 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_6 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_6 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_6 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_6 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_6 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_6 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_6 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_6 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_6 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_6 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_6 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_6 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_6 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_6 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_6 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_6 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_6 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_6 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_6 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_6 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_6 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_6 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_6 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_6 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_6 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_6 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_6 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_6 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_6 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_6 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_6 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_6 = invSboxRom_254;
      default : _zz__zz_stateReg_75_6 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_9)
      8'b00000000 : _zz__zz_stateReg_75_8 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_8 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_8 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_8 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_8 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_8 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_8 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_8 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_8 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_8 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_8 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_8 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_8 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_8 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_8 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_8 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_8 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_8 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_8 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_8 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_8 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_8 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_8 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_8 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_8 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_8 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_8 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_8 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_8 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_8 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_8 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_8 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_8 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_8 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_8 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_8 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_8 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_8 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_8 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_8 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_8 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_8 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_8 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_8 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_8 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_8 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_8 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_8 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_8 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_8 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_8 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_8 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_8 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_8 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_8 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_8 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_8 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_8 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_8 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_8 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_8 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_8 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_8 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_8 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_8 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_8 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_8 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_8 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_8 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_8 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_8 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_8 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_8 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_8 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_8 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_8 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_8 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_8 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_8 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_8 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_8 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_8 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_8 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_8 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_8 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_8 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_8 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_8 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_8 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_8 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_8 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_8 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_8 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_8 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_8 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_8 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_8 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_8 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_8 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_8 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_8 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_8 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_8 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_8 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_8 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_8 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_8 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_8 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_8 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_8 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_8 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_8 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_8 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_8 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_8 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_8 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_8 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_8 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_8 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_8 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_8 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_8 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_8 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_8 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_8 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_8 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_8 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_8 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_8 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_8 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_8 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_8 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_8 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_8 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_8 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_8 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_8 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_8 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_8 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_8 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_8 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_8 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_8 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_8 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_8 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_8 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_8 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_8 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_8 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_8 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_8 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_8 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_8 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_8 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_8 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_8 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_8 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_8 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_8 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_8 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_8 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_8 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_8 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_8 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_8 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_8 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_8 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_8 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_8 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_8 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_8 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_8 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_8 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_8 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_8 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_8 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_8 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_8 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_8 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_8 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_8 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_8 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_8 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_8 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_8 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_8 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_8 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_8 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_8 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_8 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_8 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_8 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_8 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_8 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_8 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_8 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_8 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_8 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_8 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_8 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_8 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_8 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_8 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_8 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_8 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_8 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_8 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_8 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_8 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_8 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_8 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_8 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_8 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_8 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_8 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_8 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_8 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_8 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_8 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_8 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_8 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_8 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_8 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_8 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_8 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_8 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_8 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_8 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_8 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_8 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_8 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_8 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_8 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_8 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_8 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_8 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_8 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_8 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_8 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_8 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_8 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_8 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_8 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_8 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_8 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_8 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_8 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_8 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_8 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_8 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_8 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_8 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_8 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_8 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_8 = invSboxRom_254;
      default : _zz__zz_stateReg_75_8 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_12)
      8'b00000000 : _zz__zz_stateReg_75_11 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_11 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_11 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_11 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_11 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_11 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_11 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_11 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_11 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_11 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_11 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_11 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_11 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_11 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_11 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_11 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_11 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_11 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_11 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_11 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_11 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_11 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_11 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_11 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_11 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_11 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_11 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_11 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_11 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_11 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_11 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_11 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_11 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_11 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_11 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_11 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_11 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_11 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_11 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_11 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_11 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_11 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_11 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_11 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_11 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_11 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_11 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_11 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_11 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_11 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_11 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_11 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_11 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_11 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_11 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_11 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_11 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_11 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_11 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_11 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_11 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_11 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_11 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_11 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_11 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_11 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_11 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_11 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_11 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_11 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_11 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_11 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_11 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_11 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_11 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_11 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_11 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_11 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_11 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_11 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_11 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_11 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_11 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_11 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_11 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_11 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_11 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_11 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_11 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_11 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_11 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_11 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_11 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_11 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_11 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_11 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_11 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_11 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_11 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_11 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_11 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_11 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_11 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_11 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_11 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_11 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_11 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_11 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_11 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_11 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_11 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_11 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_11 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_11 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_11 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_11 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_11 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_11 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_11 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_11 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_11 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_11 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_11 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_11 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_11 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_11 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_11 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_11 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_11 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_11 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_11 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_11 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_11 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_11 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_11 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_11 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_11 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_11 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_11 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_11 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_11 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_11 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_11 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_11 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_11 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_11 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_11 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_11 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_11 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_11 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_11 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_11 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_11 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_11 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_11 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_11 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_11 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_11 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_11 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_11 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_11 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_11 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_11 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_11 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_11 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_11 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_11 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_11 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_11 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_11 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_11 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_11 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_11 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_11 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_11 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_11 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_11 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_11 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_11 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_11 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_11 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_11 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_11 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_11 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_11 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_11 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_11 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_11 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_11 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_11 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_11 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_11 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_11 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_11 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_11 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_11 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_11 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_11 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_11 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_11 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_11 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_11 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_11 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_11 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_11 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_11 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_11 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_11 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_11 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_11 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_11 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_11 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_11 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_11 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_11 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_11 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_11 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_11 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_11 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_11 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_11 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_11 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_11 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_11 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_11 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_11 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_11 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_11 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_11 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_11 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_11 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_11 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_11 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_11 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_11 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_11 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_11 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_11 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_11 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_11 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_11 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_11 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_11 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_11 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_11 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_11 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_11 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_11 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_11 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_11 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_11 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_11 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_11 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_11 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_11 = invSboxRom_254;
      default : _zz__zz_stateReg_75_11 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_14)
      8'b00000000 : _zz__zz_stateReg_75_13 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_13 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_13 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_13 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_13 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_13 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_13 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_13 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_13 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_13 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_13 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_13 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_13 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_13 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_13 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_13 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_13 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_13 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_13 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_13 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_13 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_13 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_13 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_13 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_13 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_13 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_13 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_13 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_13 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_13 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_13 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_13 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_13 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_13 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_13 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_13 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_13 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_13 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_13 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_13 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_13 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_13 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_13 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_13 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_13 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_13 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_13 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_13 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_13 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_13 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_13 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_13 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_13 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_13 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_13 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_13 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_13 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_13 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_13 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_13 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_13 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_13 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_13 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_13 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_13 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_13 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_13 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_13 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_13 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_13 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_13 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_13 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_13 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_13 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_13 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_13 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_13 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_13 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_13 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_13 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_13 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_13 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_13 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_13 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_13 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_13 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_13 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_13 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_13 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_13 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_13 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_13 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_13 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_13 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_13 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_13 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_13 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_13 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_13 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_13 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_13 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_13 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_13 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_13 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_13 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_13 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_13 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_13 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_13 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_13 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_13 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_13 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_13 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_13 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_13 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_13 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_13 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_13 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_13 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_13 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_13 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_13 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_13 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_13 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_13 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_13 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_13 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_13 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_13 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_13 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_13 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_13 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_13 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_13 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_13 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_13 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_13 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_13 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_13 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_13 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_13 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_13 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_13 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_13 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_13 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_13 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_13 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_13 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_13 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_13 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_13 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_13 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_13 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_13 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_13 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_13 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_13 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_13 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_13 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_13 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_13 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_13 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_13 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_13 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_13 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_13 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_13 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_13 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_13 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_13 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_13 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_13 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_13 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_13 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_13 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_13 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_13 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_13 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_13 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_13 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_13 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_13 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_13 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_13 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_13 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_13 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_13 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_13 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_13 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_13 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_13 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_13 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_13 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_13 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_13 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_13 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_13 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_13 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_13 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_13 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_13 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_13 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_13 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_13 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_13 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_13 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_13 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_13 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_13 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_13 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_13 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_13 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_13 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_13 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_13 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_13 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_13 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_13 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_13 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_13 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_13 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_13 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_13 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_13 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_13 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_13 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_13 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_13 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_13 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_13 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_13 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_13 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_13 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_13 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_13 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_13 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_13 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_13 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_13 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_13 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_13 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_13 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_13 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_13 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_13 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_13 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_13 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_13 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_13 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_13 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_13 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_13 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_13 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_13 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_13 = invSboxRom_254;
      default : _zz__zz_stateReg_75_13 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_16)
      8'b00000000 : _zz__zz_stateReg_75_15 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_15 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_15 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_15 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_15 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_15 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_15 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_15 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_15 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_15 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_15 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_15 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_15 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_15 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_15 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_15 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_15 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_15 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_15 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_15 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_15 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_15 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_15 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_15 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_15 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_15 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_15 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_15 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_15 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_15 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_15 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_15 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_15 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_15 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_15 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_15 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_15 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_15 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_15 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_15 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_15 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_15 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_15 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_15 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_15 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_15 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_15 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_15 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_15 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_15 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_15 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_15 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_15 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_15 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_15 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_15 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_15 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_15 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_15 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_15 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_15 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_15 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_15 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_15 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_15 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_15 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_15 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_15 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_15 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_15 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_15 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_15 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_15 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_15 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_15 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_15 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_15 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_15 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_15 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_15 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_15 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_15 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_15 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_15 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_15 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_15 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_15 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_15 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_15 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_15 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_15 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_15 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_15 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_15 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_15 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_15 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_15 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_15 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_15 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_15 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_15 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_15 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_15 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_15 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_15 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_15 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_15 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_15 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_15 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_15 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_15 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_15 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_15 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_15 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_15 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_15 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_15 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_15 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_15 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_15 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_15 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_15 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_15 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_15 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_15 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_15 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_15 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_15 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_15 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_15 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_15 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_15 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_15 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_15 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_15 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_15 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_15 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_15 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_15 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_15 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_15 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_15 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_15 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_15 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_15 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_15 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_15 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_15 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_15 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_15 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_15 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_15 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_15 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_15 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_15 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_15 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_15 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_15 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_15 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_15 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_15 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_15 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_15 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_15 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_15 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_15 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_15 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_15 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_15 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_15 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_15 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_15 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_15 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_15 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_15 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_15 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_15 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_15 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_15 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_15 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_15 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_15 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_15 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_15 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_15 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_15 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_15 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_15 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_15 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_15 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_15 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_15 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_15 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_15 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_15 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_15 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_15 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_15 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_15 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_15 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_15 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_15 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_15 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_15 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_15 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_15 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_15 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_15 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_15 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_15 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_15 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_15 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_15 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_15 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_15 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_15 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_15 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_15 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_15 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_15 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_15 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_15 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_15 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_15 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_15 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_15 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_15 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_15 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_15 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_15 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_15 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_15 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_15 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_15 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_15 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_15 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_15 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_15 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_15 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_15 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_15 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_15 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_15 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_15 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_15 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_15 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_15 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_15 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_15 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_15 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_15 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_15 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_15 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_15 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_15 = invSboxRom_254;
      default : _zz__zz_stateReg_75_15 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_18)
      8'b00000000 : _zz__zz_stateReg_75_17 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_17 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_17 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_17 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_17 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_17 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_17 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_17 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_17 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_17 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_17 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_17 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_17 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_17 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_17 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_17 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_17 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_17 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_17 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_17 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_17 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_17 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_17 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_17 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_17 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_17 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_17 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_17 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_17 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_17 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_17 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_17 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_17 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_17 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_17 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_17 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_17 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_17 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_17 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_17 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_17 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_17 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_17 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_17 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_17 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_17 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_17 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_17 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_17 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_17 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_17 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_17 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_17 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_17 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_17 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_17 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_17 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_17 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_17 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_17 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_17 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_17 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_17 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_17 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_17 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_17 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_17 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_17 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_17 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_17 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_17 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_17 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_17 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_17 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_17 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_17 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_17 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_17 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_17 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_17 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_17 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_17 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_17 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_17 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_17 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_17 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_17 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_17 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_17 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_17 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_17 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_17 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_17 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_17 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_17 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_17 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_17 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_17 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_17 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_17 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_17 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_17 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_17 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_17 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_17 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_17 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_17 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_17 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_17 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_17 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_17 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_17 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_17 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_17 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_17 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_17 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_17 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_17 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_17 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_17 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_17 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_17 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_17 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_17 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_17 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_17 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_17 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_17 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_17 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_17 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_17 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_17 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_17 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_17 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_17 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_17 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_17 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_17 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_17 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_17 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_17 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_17 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_17 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_17 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_17 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_17 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_17 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_17 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_17 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_17 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_17 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_17 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_17 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_17 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_17 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_17 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_17 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_17 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_17 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_17 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_17 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_17 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_17 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_17 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_17 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_17 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_17 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_17 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_17 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_17 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_17 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_17 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_17 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_17 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_17 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_17 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_17 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_17 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_17 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_17 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_17 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_17 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_17 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_17 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_17 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_17 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_17 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_17 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_17 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_17 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_17 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_17 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_17 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_17 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_17 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_17 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_17 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_17 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_17 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_17 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_17 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_17 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_17 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_17 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_17 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_17 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_17 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_17 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_17 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_17 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_17 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_17 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_17 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_17 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_17 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_17 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_17 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_17 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_17 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_17 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_17 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_17 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_17 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_17 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_17 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_17 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_17 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_17 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_17 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_17 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_17 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_17 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_17 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_17 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_17 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_17 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_17 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_17 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_17 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_17 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_17 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_17 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_17 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_17 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_17 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_17 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_17 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_17 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_17 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_17 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_17 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_17 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_17 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_17 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_17 = invSboxRom_254;
      default : _zz__zz_stateReg_75_17 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_20)
      8'b00000000 : _zz__zz_stateReg_75_19 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_19 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_19 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_19 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_19 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_19 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_19 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_19 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_19 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_19 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_19 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_19 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_19 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_19 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_19 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_19 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_19 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_19 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_19 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_19 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_19 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_19 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_19 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_19 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_19 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_19 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_19 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_19 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_19 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_19 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_19 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_19 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_19 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_19 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_19 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_19 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_19 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_19 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_19 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_19 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_19 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_19 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_19 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_19 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_19 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_19 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_19 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_19 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_19 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_19 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_19 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_19 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_19 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_19 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_19 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_19 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_19 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_19 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_19 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_19 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_19 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_19 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_19 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_19 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_19 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_19 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_19 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_19 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_19 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_19 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_19 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_19 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_19 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_19 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_19 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_19 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_19 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_19 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_19 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_19 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_19 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_19 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_19 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_19 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_19 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_19 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_19 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_19 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_19 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_19 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_19 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_19 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_19 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_19 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_19 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_19 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_19 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_19 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_19 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_19 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_19 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_19 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_19 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_19 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_19 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_19 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_19 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_19 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_19 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_19 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_19 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_19 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_19 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_19 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_19 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_19 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_19 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_19 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_19 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_19 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_19 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_19 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_19 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_19 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_19 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_19 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_19 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_19 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_19 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_19 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_19 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_19 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_19 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_19 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_19 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_19 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_19 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_19 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_19 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_19 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_19 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_19 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_19 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_19 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_19 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_19 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_19 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_19 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_19 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_19 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_19 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_19 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_19 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_19 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_19 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_19 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_19 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_19 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_19 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_19 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_19 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_19 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_19 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_19 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_19 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_19 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_19 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_19 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_19 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_19 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_19 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_19 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_19 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_19 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_19 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_19 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_19 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_19 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_19 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_19 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_19 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_19 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_19 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_19 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_19 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_19 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_19 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_19 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_19 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_19 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_19 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_19 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_19 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_19 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_19 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_19 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_19 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_19 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_19 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_19 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_19 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_19 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_19 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_19 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_19 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_19 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_19 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_19 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_19 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_19 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_19 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_19 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_19 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_19 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_19 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_19 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_19 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_19 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_19 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_19 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_19 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_19 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_19 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_19 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_19 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_19 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_19 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_19 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_19 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_19 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_19 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_19 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_19 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_19 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_19 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_19 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_19 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_19 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_19 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_19 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_19 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_19 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_19 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_19 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_19 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_19 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_19 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_19 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_19 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_19 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_19 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_19 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_19 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_19 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_19 = invSboxRom_254;
      default : _zz__zz_stateReg_75_19 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_22)
      8'b00000000 : _zz__zz_stateReg_75_21 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_21 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_21 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_21 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_21 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_21 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_21 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_21 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_21 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_21 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_21 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_21 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_21 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_21 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_21 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_21 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_21 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_21 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_21 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_21 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_21 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_21 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_21 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_21 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_21 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_21 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_21 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_21 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_21 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_21 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_21 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_21 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_21 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_21 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_21 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_21 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_21 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_21 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_21 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_21 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_21 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_21 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_21 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_21 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_21 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_21 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_21 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_21 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_21 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_21 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_21 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_21 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_21 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_21 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_21 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_21 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_21 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_21 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_21 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_21 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_21 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_21 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_21 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_21 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_21 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_21 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_21 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_21 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_21 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_21 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_21 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_21 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_21 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_21 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_21 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_21 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_21 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_21 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_21 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_21 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_21 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_21 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_21 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_21 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_21 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_21 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_21 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_21 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_21 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_21 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_21 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_21 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_21 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_21 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_21 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_21 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_21 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_21 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_21 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_21 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_21 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_21 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_21 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_21 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_21 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_21 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_21 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_21 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_21 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_21 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_21 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_21 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_21 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_21 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_21 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_21 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_21 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_21 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_21 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_21 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_21 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_21 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_21 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_21 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_21 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_21 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_21 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_21 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_21 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_21 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_21 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_21 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_21 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_21 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_21 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_21 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_21 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_21 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_21 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_21 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_21 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_21 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_21 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_21 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_21 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_21 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_21 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_21 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_21 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_21 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_21 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_21 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_21 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_21 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_21 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_21 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_21 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_21 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_21 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_21 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_21 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_21 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_21 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_21 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_21 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_21 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_21 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_21 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_21 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_21 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_21 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_21 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_21 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_21 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_21 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_21 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_21 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_21 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_21 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_21 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_21 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_21 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_21 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_21 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_21 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_21 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_21 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_21 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_21 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_21 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_21 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_21 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_21 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_21 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_21 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_21 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_21 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_21 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_21 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_21 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_21 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_21 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_21 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_21 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_21 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_21 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_21 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_21 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_21 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_21 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_21 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_21 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_21 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_21 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_21 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_21 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_21 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_21 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_21 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_21 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_21 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_21 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_21 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_21 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_21 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_21 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_21 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_21 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_21 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_21 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_21 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_21 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_21 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_21 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_21 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_21 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_21 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_21 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_21 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_21 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_21 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_21 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_21 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_21 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_21 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_21 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_21 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_21 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_21 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_21 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_21 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_21 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_21 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_21 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_21 = invSboxRom_254;
      default : _zz__zz_stateReg_75_21 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_25)
      8'b00000000 : _zz__zz_stateReg_75_24 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_24 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_24 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_24 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_24 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_24 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_24 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_24 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_24 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_24 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_24 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_24 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_24 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_24 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_24 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_24 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_24 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_24 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_24 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_24 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_24 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_24 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_24 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_24 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_24 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_24 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_24 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_24 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_24 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_24 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_24 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_24 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_24 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_24 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_24 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_24 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_24 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_24 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_24 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_24 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_24 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_24 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_24 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_24 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_24 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_24 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_24 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_24 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_24 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_24 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_24 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_24 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_24 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_24 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_24 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_24 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_24 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_24 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_24 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_24 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_24 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_24 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_24 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_24 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_24 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_24 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_24 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_24 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_24 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_24 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_24 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_24 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_24 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_24 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_24 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_24 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_24 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_24 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_24 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_24 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_24 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_24 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_24 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_24 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_24 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_24 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_24 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_24 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_24 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_24 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_24 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_24 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_24 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_24 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_24 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_24 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_24 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_24 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_24 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_24 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_24 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_24 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_24 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_24 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_24 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_24 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_24 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_24 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_24 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_24 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_24 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_24 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_24 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_24 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_24 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_24 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_24 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_24 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_24 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_24 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_24 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_24 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_24 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_24 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_24 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_24 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_24 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_24 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_24 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_24 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_24 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_24 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_24 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_24 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_24 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_24 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_24 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_24 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_24 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_24 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_24 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_24 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_24 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_24 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_24 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_24 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_24 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_24 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_24 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_24 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_24 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_24 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_24 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_24 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_24 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_24 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_24 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_24 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_24 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_24 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_24 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_24 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_24 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_24 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_24 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_24 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_24 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_24 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_24 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_24 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_24 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_24 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_24 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_24 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_24 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_24 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_24 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_24 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_24 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_24 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_24 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_24 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_24 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_24 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_24 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_24 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_24 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_24 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_24 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_24 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_24 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_24 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_24 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_24 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_24 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_24 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_24 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_24 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_24 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_24 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_24 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_24 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_24 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_24 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_24 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_24 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_24 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_24 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_24 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_24 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_24 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_24 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_24 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_24 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_24 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_24 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_24 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_24 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_24 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_24 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_24 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_24 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_24 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_24 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_24 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_24 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_24 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_24 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_24 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_24 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_24 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_24 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_24 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_24 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_24 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_24 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_24 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_24 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_24 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_24 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_24 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_24 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_24 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_24 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_24 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_24 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_24 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_24 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_24 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_24 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_24 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_24 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_24 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_24 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_24 = invSboxRom_254;
      default : _zz__zz_stateReg_75_24 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_27)
      8'b00000000 : _zz__zz_stateReg_75_26 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_26 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_26 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_26 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_26 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_26 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_26 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_26 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_26 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_26 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_26 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_26 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_26 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_26 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_26 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_26 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_26 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_26 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_26 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_26 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_26 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_26 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_26 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_26 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_26 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_26 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_26 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_26 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_26 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_26 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_26 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_26 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_26 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_26 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_26 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_26 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_26 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_26 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_26 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_26 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_26 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_26 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_26 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_26 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_26 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_26 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_26 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_26 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_26 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_26 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_26 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_26 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_26 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_26 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_26 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_26 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_26 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_26 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_26 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_26 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_26 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_26 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_26 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_26 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_26 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_26 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_26 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_26 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_26 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_26 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_26 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_26 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_26 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_26 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_26 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_26 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_26 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_26 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_26 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_26 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_26 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_26 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_26 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_26 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_26 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_26 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_26 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_26 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_26 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_26 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_26 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_26 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_26 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_26 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_26 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_26 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_26 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_26 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_26 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_26 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_26 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_26 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_26 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_26 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_26 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_26 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_26 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_26 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_26 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_26 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_26 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_26 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_26 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_26 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_26 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_26 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_26 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_26 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_26 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_26 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_26 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_26 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_26 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_26 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_26 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_26 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_26 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_26 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_26 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_26 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_26 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_26 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_26 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_26 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_26 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_26 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_26 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_26 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_26 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_26 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_26 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_26 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_26 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_26 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_26 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_26 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_26 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_26 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_26 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_26 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_26 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_26 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_26 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_26 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_26 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_26 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_26 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_26 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_26 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_26 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_26 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_26 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_26 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_26 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_26 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_26 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_26 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_26 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_26 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_26 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_26 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_26 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_26 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_26 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_26 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_26 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_26 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_26 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_26 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_26 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_26 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_26 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_26 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_26 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_26 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_26 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_26 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_26 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_26 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_26 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_26 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_26 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_26 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_26 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_26 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_26 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_26 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_26 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_26 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_26 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_26 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_26 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_26 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_26 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_26 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_26 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_26 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_26 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_26 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_26 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_26 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_26 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_26 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_26 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_26 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_26 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_26 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_26 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_26 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_26 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_26 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_26 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_26 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_26 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_26 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_26 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_26 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_26 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_26 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_26 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_26 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_26 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_26 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_26 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_26 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_26 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_26 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_26 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_26 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_26 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_26 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_26 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_26 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_26 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_26 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_26 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_26 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_26 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_26 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_26 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_26 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_26 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_26 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_26 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_26 = invSboxRom_254;
      default : _zz__zz_stateReg_75_26 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_29)
      8'b00000000 : _zz__zz_stateReg_75_28 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_28 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_28 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_28 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_28 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_28 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_28 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_28 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_28 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_28 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_28 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_28 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_28 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_28 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_28 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_28 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_28 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_28 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_28 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_28 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_28 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_28 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_28 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_28 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_28 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_28 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_28 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_28 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_28 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_28 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_28 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_28 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_28 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_28 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_28 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_28 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_28 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_28 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_28 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_28 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_28 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_28 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_28 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_28 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_28 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_28 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_28 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_28 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_28 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_28 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_28 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_28 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_28 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_28 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_28 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_28 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_28 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_28 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_28 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_28 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_28 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_28 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_28 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_28 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_28 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_28 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_28 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_28 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_28 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_28 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_28 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_28 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_28 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_28 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_28 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_28 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_28 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_28 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_28 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_28 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_28 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_28 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_28 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_28 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_28 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_28 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_28 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_28 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_28 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_28 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_28 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_28 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_28 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_28 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_28 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_28 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_28 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_28 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_28 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_28 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_28 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_28 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_28 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_28 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_28 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_28 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_28 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_28 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_28 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_28 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_28 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_28 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_28 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_28 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_28 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_28 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_28 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_28 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_28 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_28 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_28 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_28 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_28 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_28 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_28 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_28 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_28 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_28 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_28 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_28 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_28 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_28 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_28 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_28 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_28 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_28 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_28 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_28 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_28 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_28 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_28 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_28 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_28 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_28 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_28 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_28 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_28 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_28 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_28 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_28 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_28 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_28 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_28 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_28 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_28 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_28 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_28 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_28 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_28 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_28 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_28 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_28 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_28 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_28 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_28 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_28 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_28 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_28 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_28 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_28 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_28 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_28 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_28 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_28 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_28 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_28 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_28 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_28 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_28 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_28 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_28 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_28 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_28 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_28 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_28 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_28 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_28 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_28 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_28 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_28 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_28 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_28 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_28 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_28 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_28 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_28 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_28 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_28 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_28 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_28 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_28 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_28 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_28 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_28 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_28 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_28 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_28 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_28 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_28 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_28 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_28 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_28 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_28 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_28 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_28 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_28 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_28 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_28 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_28 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_28 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_28 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_28 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_28 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_28 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_28 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_28 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_28 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_28 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_28 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_28 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_28 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_28 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_28 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_28 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_28 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_28 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_28 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_28 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_28 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_28 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_28 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_28 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_28 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_28 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_28 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_28 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_28 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_28 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_28 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_28 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_28 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_28 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_28 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_28 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_28 = invSboxRom_254;
      default : _zz__zz_stateReg_75_28 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_31)
      8'b00000000 : _zz__zz_stateReg_75_30 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_30 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_30 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_30 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_30 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_30 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_30 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_30 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_30 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_30 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_30 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_30 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_30 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_30 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_30 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_30 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_30 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_30 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_30 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_30 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_30 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_30 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_30 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_30 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_30 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_30 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_30 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_30 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_30 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_30 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_30 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_30 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_30 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_30 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_30 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_30 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_30 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_30 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_30 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_30 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_30 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_30 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_30 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_30 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_30 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_30 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_30 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_30 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_30 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_30 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_30 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_30 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_30 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_30 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_30 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_30 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_30 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_30 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_30 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_30 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_30 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_30 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_30 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_30 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_30 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_30 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_30 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_30 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_30 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_30 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_30 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_30 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_30 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_30 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_30 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_30 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_30 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_30 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_30 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_30 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_30 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_30 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_30 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_30 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_30 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_30 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_30 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_30 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_30 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_30 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_30 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_30 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_30 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_30 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_30 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_30 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_30 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_30 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_30 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_30 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_30 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_30 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_30 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_30 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_30 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_30 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_30 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_30 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_30 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_30 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_30 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_30 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_30 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_30 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_30 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_30 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_30 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_30 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_30 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_30 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_30 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_30 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_30 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_30 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_30 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_30 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_30 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_30 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_30 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_30 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_30 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_30 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_30 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_30 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_30 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_30 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_30 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_30 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_30 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_30 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_30 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_30 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_30 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_30 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_30 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_30 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_30 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_30 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_30 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_30 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_30 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_30 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_30 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_30 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_30 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_30 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_30 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_30 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_30 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_30 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_30 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_30 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_30 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_30 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_30 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_30 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_30 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_30 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_30 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_30 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_30 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_30 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_30 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_30 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_30 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_30 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_30 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_30 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_30 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_30 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_30 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_30 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_30 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_30 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_30 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_30 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_30 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_30 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_30 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_30 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_30 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_30 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_30 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_30 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_30 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_30 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_30 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_30 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_30 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_30 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_30 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_30 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_30 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_30 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_30 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_30 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_30 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_30 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_30 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_30 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_30 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_30 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_30 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_30 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_30 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_30 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_30 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_30 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_30 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_30 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_30 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_30 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_30 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_30 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_30 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_30 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_30 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_30 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_30 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_30 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_30 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_30 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_30 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_30 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_30 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_30 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_30 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_30 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_30 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_30 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_30 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_30 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_30 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_30 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_30 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_30 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_30 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_30 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_30 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_30 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_30 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_30 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_30 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_30 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_30 = invSboxRom_254;
      default : _zz__zz_stateReg_75_30 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_33)
      8'b00000000 : _zz__zz_stateReg_75_32 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_32 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_32 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_32 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_32 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_32 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_32 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_32 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_32 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_32 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_32 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_32 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_32 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_32 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_32 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_32 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_32 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_32 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_32 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_32 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_32 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_32 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_32 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_32 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_32 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_32 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_32 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_32 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_32 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_32 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_32 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_32 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_32 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_32 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_32 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_32 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_32 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_32 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_32 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_32 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_32 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_32 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_32 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_32 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_32 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_32 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_32 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_32 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_32 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_32 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_32 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_32 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_32 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_32 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_32 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_32 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_32 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_32 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_32 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_32 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_32 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_32 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_32 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_32 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_32 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_32 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_32 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_32 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_32 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_32 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_32 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_32 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_32 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_32 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_32 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_32 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_32 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_32 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_32 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_32 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_32 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_32 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_32 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_32 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_32 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_32 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_32 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_32 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_32 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_32 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_32 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_32 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_32 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_32 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_32 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_32 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_32 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_32 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_32 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_32 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_32 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_32 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_32 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_32 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_32 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_32 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_32 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_32 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_32 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_32 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_32 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_32 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_32 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_32 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_32 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_32 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_32 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_32 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_32 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_32 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_32 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_32 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_32 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_32 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_32 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_32 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_32 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_32 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_32 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_32 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_32 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_32 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_32 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_32 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_32 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_32 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_32 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_32 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_32 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_32 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_32 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_32 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_32 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_32 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_32 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_32 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_32 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_32 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_32 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_32 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_32 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_32 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_32 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_32 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_32 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_32 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_32 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_32 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_32 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_32 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_32 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_32 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_32 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_32 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_32 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_32 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_32 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_32 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_32 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_32 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_32 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_32 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_32 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_32 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_32 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_32 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_32 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_32 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_32 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_32 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_32 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_32 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_32 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_32 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_32 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_32 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_32 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_32 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_32 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_32 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_32 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_32 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_32 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_32 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_32 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_32 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_32 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_32 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_32 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_32 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_32 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_32 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_32 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_32 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_32 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_32 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_32 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_32 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_32 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_32 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_32 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_32 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_32 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_32 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_32 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_32 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_32 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_32 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_32 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_32 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_32 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_32 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_32 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_32 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_32 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_32 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_32 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_32 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_32 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_32 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_32 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_32 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_32 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_32 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_32 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_32 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_32 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_32 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_32 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_32 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_32 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_32 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_32 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_32 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_32 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_32 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_32 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_32 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_32 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_32 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_32 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_32 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_32 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_32 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_32 = invSboxRom_254;
      default : _zz__zz_stateReg_75_32 = invSboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_75_35)
      8'b00000000 : _zz__zz_stateReg_75_34 = invSboxRom_0;
      8'b00000001 : _zz__zz_stateReg_75_34 = invSboxRom_1;
      8'b00000010 : _zz__zz_stateReg_75_34 = invSboxRom_2;
      8'b00000011 : _zz__zz_stateReg_75_34 = invSboxRom_3;
      8'b00000100 : _zz__zz_stateReg_75_34 = invSboxRom_4;
      8'b00000101 : _zz__zz_stateReg_75_34 = invSboxRom_5;
      8'b00000110 : _zz__zz_stateReg_75_34 = invSboxRom_6;
      8'b00000111 : _zz__zz_stateReg_75_34 = invSboxRom_7;
      8'b00001000 : _zz__zz_stateReg_75_34 = invSboxRom_8;
      8'b00001001 : _zz__zz_stateReg_75_34 = invSboxRom_9;
      8'b00001010 : _zz__zz_stateReg_75_34 = invSboxRom_10;
      8'b00001011 : _zz__zz_stateReg_75_34 = invSboxRom_11;
      8'b00001100 : _zz__zz_stateReg_75_34 = invSboxRom_12;
      8'b00001101 : _zz__zz_stateReg_75_34 = invSboxRom_13;
      8'b00001110 : _zz__zz_stateReg_75_34 = invSboxRom_14;
      8'b00001111 : _zz__zz_stateReg_75_34 = invSboxRom_15;
      8'b00010000 : _zz__zz_stateReg_75_34 = invSboxRom_16;
      8'b00010001 : _zz__zz_stateReg_75_34 = invSboxRom_17;
      8'b00010010 : _zz__zz_stateReg_75_34 = invSboxRom_18;
      8'b00010011 : _zz__zz_stateReg_75_34 = invSboxRom_19;
      8'b00010100 : _zz__zz_stateReg_75_34 = invSboxRom_20;
      8'b00010101 : _zz__zz_stateReg_75_34 = invSboxRom_21;
      8'b00010110 : _zz__zz_stateReg_75_34 = invSboxRom_22;
      8'b00010111 : _zz__zz_stateReg_75_34 = invSboxRom_23;
      8'b00011000 : _zz__zz_stateReg_75_34 = invSboxRom_24;
      8'b00011001 : _zz__zz_stateReg_75_34 = invSboxRom_25;
      8'b00011010 : _zz__zz_stateReg_75_34 = invSboxRom_26;
      8'b00011011 : _zz__zz_stateReg_75_34 = invSboxRom_27;
      8'b00011100 : _zz__zz_stateReg_75_34 = invSboxRom_28;
      8'b00011101 : _zz__zz_stateReg_75_34 = invSboxRom_29;
      8'b00011110 : _zz__zz_stateReg_75_34 = invSboxRom_30;
      8'b00011111 : _zz__zz_stateReg_75_34 = invSboxRom_31;
      8'b00100000 : _zz__zz_stateReg_75_34 = invSboxRom_32;
      8'b00100001 : _zz__zz_stateReg_75_34 = invSboxRom_33;
      8'b00100010 : _zz__zz_stateReg_75_34 = invSboxRom_34;
      8'b00100011 : _zz__zz_stateReg_75_34 = invSboxRom_35;
      8'b00100100 : _zz__zz_stateReg_75_34 = invSboxRom_36;
      8'b00100101 : _zz__zz_stateReg_75_34 = invSboxRom_37;
      8'b00100110 : _zz__zz_stateReg_75_34 = invSboxRom_38;
      8'b00100111 : _zz__zz_stateReg_75_34 = invSboxRom_39;
      8'b00101000 : _zz__zz_stateReg_75_34 = invSboxRom_40;
      8'b00101001 : _zz__zz_stateReg_75_34 = invSboxRom_41;
      8'b00101010 : _zz__zz_stateReg_75_34 = invSboxRom_42;
      8'b00101011 : _zz__zz_stateReg_75_34 = invSboxRom_43;
      8'b00101100 : _zz__zz_stateReg_75_34 = invSboxRom_44;
      8'b00101101 : _zz__zz_stateReg_75_34 = invSboxRom_45;
      8'b00101110 : _zz__zz_stateReg_75_34 = invSboxRom_46;
      8'b00101111 : _zz__zz_stateReg_75_34 = invSboxRom_47;
      8'b00110000 : _zz__zz_stateReg_75_34 = invSboxRom_48;
      8'b00110001 : _zz__zz_stateReg_75_34 = invSboxRom_49;
      8'b00110010 : _zz__zz_stateReg_75_34 = invSboxRom_50;
      8'b00110011 : _zz__zz_stateReg_75_34 = invSboxRom_51;
      8'b00110100 : _zz__zz_stateReg_75_34 = invSboxRom_52;
      8'b00110101 : _zz__zz_stateReg_75_34 = invSboxRom_53;
      8'b00110110 : _zz__zz_stateReg_75_34 = invSboxRom_54;
      8'b00110111 : _zz__zz_stateReg_75_34 = invSboxRom_55;
      8'b00111000 : _zz__zz_stateReg_75_34 = invSboxRom_56;
      8'b00111001 : _zz__zz_stateReg_75_34 = invSboxRom_57;
      8'b00111010 : _zz__zz_stateReg_75_34 = invSboxRom_58;
      8'b00111011 : _zz__zz_stateReg_75_34 = invSboxRom_59;
      8'b00111100 : _zz__zz_stateReg_75_34 = invSboxRom_60;
      8'b00111101 : _zz__zz_stateReg_75_34 = invSboxRom_61;
      8'b00111110 : _zz__zz_stateReg_75_34 = invSboxRom_62;
      8'b00111111 : _zz__zz_stateReg_75_34 = invSboxRom_63;
      8'b01000000 : _zz__zz_stateReg_75_34 = invSboxRom_64;
      8'b01000001 : _zz__zz_stateReg_75_34 = invSboxRom_65;
      8'b01000010 : _zz__zz_stateReg_75_34 = invSboxRom_66;
      8'b01000011 : _zz__zz_stateReg_75_34 = invSboxRom_67;
      8'b01000100 : _zz__zz_stateReg_75_34 = invSboxRom_68;
      8'b01000101 : _zz__zz_stateReg_75_34 = invSboxRom_69;
      8'b01000110 : _zz__zz_stateReg_75_34 = invSboxRom_70;
      8'b01000111 : _zz__zz_stateReg_75_34 = invSboxRom_71;
      8'b01001000 : _zz__zz_stateReg_75_34 = invSboxRom_72;
      8'b01001001 : _zz__zz_stateReg_75_34 = invSboxRom_73;
      8'b01001010 : _zz__zz_stateReg_75_34 = invSboxRom_74;
      8'b01001011 : _zz__zz_stateReg_75_34 = invSboxRom_75;
      8'b01001100 : _zz__zz_stateReg_75_34 = invSboxRom_76;
      8'b01001101 : _zz__zz_stateReg_75_34 = invSboxRom_77;
      8'b01001110 : _zz__zz_stateReg_75_34 = invSboxRom_78;
      8'b01001111 : _zz__zz_stateReg_75_34 = invSboxRom_79;
      8'b01010000 : _zz__zz_stateReg_75_34 = invSboxRom_80;
      8'b01010001 : _zz__zz_stateReg_75_34 = invSboxRom_81;
      8'b01010010 : _zz__zz_stateReg_75_34 = invSboxRom_82;
      8'b01010011 : _zz__zz_stateReg_75_34 = invSboxRom_83;
      8'b01010100 : _zz__zz_stateReg_75_34 = invSboxRom_84;
      8'b01010101 : _zz__zz_stateReg_75_34 = invSboxRom_85;
      8'b01010110 : _zz__zz_stateReg_75_34 = invSboxRom_86;
      8'b01010111 : _zz__zz_stateReg_75_34 = invSboxRom_87;
      8'b01011000 : _zz__zz_stateReg_75_34 = invSboxRom_88;
      8'b01011001 : _zz__zz_stateReg_75_34 = invSboxRom_89;
      8'b01011010 : _zz__zz_stateReg_75_34 = invSboxRom_90;
      8'b01011011 : _zz__zz_stateReg_75_34 = invSboxRom_91;
      8'b01011100 : _zz__zz_stateReg_75_34 = invSboxRom_92;
      8'b01011101 : _zz__zz_stateReg_75_34 = invSboxRom_93;
      8'b01011110 : _zz__zz_stateReg_75_34 = invSboxRom_94;
      8'b01011111 : _zz__zz_stateReg_75_34 = invSboxRom_95;
      8'b01100000 : _zz__zz_stateReg_75_34 = invSboxRom_96;
      8'b01100001 : _zz__zz_stateReg_75_34 = invSboxRom_97;
      8'b01100010 : _zz__zz_stateReg_75_34 = invSboxRom_98;
      8'b01100011 : _zz__zz_stateReg_75_34 = invSboxRom_99;
      8'b01100100 : _zz__zz_stateReg_75_34 = invSboxRom_100;
      8'b01100101 : _zz__zz_stateReg_75_34 = invSboxRom_101;
      8'b01100110 : _zz__zz_stateReg_75_34 = invSboxRom_102;
      8'b01100111 : _zz__zz_stateReg_75_34 = invSboxRom_103;
      8'b01101000 : _zz__zz_stateReg_75_34 = invSboxRom_104;
      8'b01101001 : _zz__zz_stateReg_75_34 = invSboxRom_105;
      8'b01101010 : _zz__zz_stateReg_75_34 = invSboxRom_106;
      8'b01101011 : _zz__zz_stateReg_75_34 = invSboxRom_107;
      8'b01101100 : _zz__zz_stateReg_75_34 = invSboxRom_108;
      8'b01101101 : _zz__zz_stateReg_75_34 = invSboxRom_109;
      8'b01101110 : _zz__zz_stateReg_75_34 = invSboxRom_110;
      8'b01101111 : _zz__zz_stateReg_75_34 = invSboxRom_111;
      8'b01110000 : _zz__zz_stateReg_75_34 = invSboxRom_112;
      8'b01110001 : _zz__zz_stateReg_75_34 = invSboxRom_113;
      8'b01110010 : _zz__zz_stateReg_75_34 = invSboxRom_114;
      8'b01110011 : _zz__zz_stateReg_75_34 = invSboxRom_115;
      8'b01110100 : _zz__zz_stateReg_75_34 = invSboxRom_116;
      8'b01110101 : _zz__zz_stateReg_75_34 = invSboxRom_117;
      8'b01110110 : _zz__zz_stateReg_75_34 = invSboxRom_118;
      8'b01110111 : _zz__zz_stateReg_75_34 = invSboxRom_119;
      8'b01111000 : _zz__zz_stateReg_75_34 = invSboxRom_120;
      8'b01111001 : _zz__zz_stateReg_75_34 = invSboxRom_121;
      8'b01111010 : _zz__zz_stateReg_75_34 = invSboxRom_122;
      8'b01111011 : _zz__zz_stateReg_75_34 = invSboxRom_123;
      8'b01111100 : _zz__zz_stateReg_75_34 = invSboxRom_124;
      8'b01111101 : _zz__zz_stateReg_75_34 = invSboxRom_125;
      8'b01111110 : _zz__zz_stateReg_75_34 = invSboxRom_126;
      8'b01111111 : _zz__zz_stateReg_75_34 = invSboxRom_127;
      8'b10000000 : _zz__zz_stateReg_75_34 = invSboxRom_128;
      8'b10000001 : _zz__zz_stateReg_75_34 = invSboxRom_129;
      8'b10000010 : _zz__zz_stateReg_75_34 = invSboxRom_130;
      8'b10000011 : _zz__zz_stateReg_75_34 = invSboxRom_131;
      8'b10000100 : _zz__zz_stateReg_75_34 = invSboxRom_132;
      8'b10000101 : _zz__zz_stateReg_75_34 = invSboxRom_133;
      8'b10000110 : _zz__zz_stateReg_75_34 = invSboxRom_134;
      8'b10000111 : _zz__zz_stateReg_75_34 = invSboxRom_135;
      8'b10001000 : _zz__zz_stateReg_75_34 = invSboxRom_136;
      8'b10001001 : _zz__zz_stateReg_75_34 = invSboxRom_137;
      8'b10001010 : _zz__zz_stateReg_75_34 = invSboxRom_138;
      8'b10001011 : _zz__zz_stateReg_75_34 = invSboxRom_139;
      8'b10001100 : _zz__zz_stateReg_75_34 = invSboxRom_140;
      8'b10001101 : _zz__zz_stateReg_75_34 = invSboxRom_141;
      8'b10001110 : _zz__zz_stateReg_75_34 = invSboxRom_142;
      8'b10001111 : _zz__zz_stateReg_75_34 = invSboxRom_143;
      8'b10010000 : _zz__zz_stateReg_75_34 = invSboxRom_144;
      8'b10010001 : _zz__zz_stateReg_75_34 = invSboxRom_145;
      8'b10010010 : _zz__zz_stateReg_75_34 = invSboxRom_146;
      8'b10010011 : _zz__zz_stateReg_75_34 = invSboxRom_147;
      8'b10010100 : _zz__zz_stateReg_75_34 = invSboxRom_148;
      8'b10010101 : _zz__zz_stateReg_75_34 = invSboxRom_149;
      8'b10010110 : _zz__zz_stateReg_75_34 = invSboxRom_150;
      8'b10010111 : _zz__zz_stateReg_75_34 = invSboxRom_151;
      8'b10011000 : _zz__zz_stateReg_75_34 = invSboxRom_152;
      8'b10011001 : _zz__zz_stateReg_75_34 = invSboxRom_153;
      8'b10011010 : _zz__zz_stateReg_75_34 = invSboxRom_154;
      8'b10011011 : _zz__zz_stateReg_75_34 = invSboxRom_155;
      8'b10011100 : _zz__zz_stateReg_75_34 = invSboxRom_156;
      8'b10011101 : _zz__zz_stateReg_75_34 = invSboxRom_157;
      8'b10011110 : _zz__zz_stateReg_75_34 = invSboxRom_158;
      8'b10011111 : _zz__zz_stateReg_75_34 = invSboxRom_159;
      8'b10100000 : _zz__zz_stateReg_75_34 = invSboxRom_160;
      8'b10100001 : _zz__zz_stateReg_75_34 = invSboxRom_161;
      8'b10100010 : _zz__zz_stateReg_75_34 = invSboxRom_162;
      8'b10100011 : _zz__zz_stateReg_75_34 = invSboxRom_163;
      8'b10100100 : _zz__zz_stateReg_75_34 = invSboxRom_164;
      8'b10100101 : _zz__zz_stateReg_75_34 = invSboxRom_165;
      8'b10100110 : _zz__zz_stateReg_75_34 = invSboxRom_166;
      8'b10100111 : _zz__zz_stateReg_75_34 = invSboxRom_167;
      8'b10101000 : _zz__zz_stateReg_75_34 = invSboxRom_168;
      8'b10101001 : _zz__zz_stateReg_75_34 = invSboxRom_169;
      8'b10101010 : _zz__zz_stateReg_75_34 = invSboxRom_170;
      8'b10101011 : _zz__zz_stateReg_75_34 = invSboxRom_171;
      8'b10101100 : _zz__zz_stateReg_75_34 = invSboxRom_172;
      8'b10101101 : _zz__zz_stateReg_75_34 = invSboxRom_173;
      8'b10101110 : _zz__zz_stateReg_75_34 = invSboxRom_174;
      8'b10101111 : _zz__zz_stateReg_75_34 = invSboxRom_175;
      8'b10110000 : _zz__zz_stateReg_75_34 = invSboxRom_176;
      8'b10110001 : _zz__zz_stateReg_75_34 = invSboxRom_177;
      8'b10110010 : _zz__zz_stateReg_75_34 = invSboxRom_178;
      8'b10110011 : _zz__zz_stateReg_75_34 = invSboxRom_179;
      8'b10110100 : _zz__zz_stateReg_75_34 = invSboxRom_180;
      8'b10110101 : _zz__zz_stateReg_75_34 = invSboxRom_181;
      8'b10110110 : _zz__zz_stateReg_75_34 = invSboxRom_182;
      8'b10110111 : _zz__zz_stateReg_75_34 = invSboxRom_183;
      8'b10111000 : _zz__zz_stateReg_75_34 = invSboxRom_184;
      8'b10111001 : _zz__zz_stateReg_75_34 = invSboxRom_185;
      8'b10111010 : _zz__zz_stateReg_75_34 = invSboxRom_186;
      8'b10111011 : _zz__zz_stateReg_75_34 = invSboxRom_187;
      8'b10111100 : _zz__zz_stateReg_75_34 = invSboxRom_188;
      8'b10111101 : _zz__zz_stateReg_75_34 = invSboxRom_189;
      8'b10111110 : _zz__zz_stateReg_75_34 = invSboxRom_190;
      8'b10111111 : _zz__zz_stateReg_75_34 = invSboxRom_191;
      8'b11000000 : _zz__zz_stateReg_75_34 = invSboxRom_192;
      8'b11000001 : _zz__zz_stateReg_75_34 = invSboxRom_193;
      8'b11000010 : _zz__zz_stateReg_75_34 = invSboxRom_194;
      8'b11000011 : _zz__zz_stateReg_75_34 = invSboxRom_195;
      8'b11000100 : _zz__zz_stateReg_75_34 = invSboxRom_196;
      8'b11000101 : _zz__zz_stateReg_75_34 = invSboxRom_197;
      8'b11000110 : _zz__zz_stateReg_75_34 = invSboxRom_198;
      8'b11000111 : _zz__zz_stateReg_75_34 = invSboxRom_199;
      8'b11001000 : _zz__zz_stateReg_75_34 = invSboxRom_200;
      8'b11001001 : _zz__zz_stateReg_75_34 = invSboxRom_201;
      8'b11001010 : _zz__zz_stateReg_75_34 = invSboxRom_202;
      8'b11001011 : _zz__zz_stateReg_75_34 = invSboxRom_203;
      8'b11001100 : _zz__zz_stateReg_75_34 = invSboxRom_204;
      8'b11001101 : _zz__zz_stateReg_75_34 = invSboxRom_205;
      8'b11001110 : _zz__zz_stateReg_75_34 = invSboxRom_206;
      8'b11001111 : _zz__zz_stateReg_75_34 = invSboxRom_207;
      8'b11010000 : _zz__zz_stateReg_75_34 = invSboxRom_208;
      8'b11010001 : _zz__zz_stateReg_75_34 = invSboxRom_209;
      8'b11010010 : _zz__zz_stateReg_75_34 = invSboxRom_210;
      8'b11010011 : _zz__zz_stateReg_75_34 = invSboxRom_211;
      8'b11010100 : _zz__zz_stateReg_75_34 = invSboxRom_212;
      8'b11010101 : _zz__zz_stateReg_75_34 = invSboxRom_213;
      8'b11010110 : _zz__zz_stateReg_75_34 = invSboxRom_214;
      8'b11010111 : _zz__zz_stateReg_75_34 = invSboxRom_215;
      8'b11011000 : _zz__zz_stateReg_75_34 = invSboxRom_216;
      8'b11011001 : _zz__zz_stateReg_75_34 = invSboxRom_217;
      8'b11011010 : _zz__zz_stateReg_75_34 = invSboxRom_218;
      8'b11011011 : _zz__zz_stateReg_75_34 = invSboxRom_219;
      8'b11011100 : _zz__zz_stateReg_75_34 = invSboxRom_220;
      8'b11011101 : _zz__zz_stateReg_75_34 = invSboxRom_221;
      8'b11011110 : _zz__zz_stateReg_75_34 = invSboxRom_222;
      8'b11011111 : _zz__zz_stateReg_75_34 = invSboxRom_223;
      8'b11100000 : _zz__zz_stateReg_75_34 = invSboxRom_224;
      8'b11100001 : _zz__zz_stateReg_75_34 = invSboxRom_225;
      8'b11100010 : _zz__zz_stateReg_75_34 = invSboxRom_226;
      8'b11100011 : _zz__zz_stateReg_75_34 = invSboxRom_227;
      8'b11100100 : _zz__zz_stateReg_75_34 = invSboxRom_228;
      8'b11100101 : _zz__zz_stateReg_75_34 = invSboxRom_229;
      8'b11100110 : _zz__zz_stateReg_75_34 = invSboxRom_230;
      8'b11100111 : _zz__zz_stateReg_75_34 = invSboxRom_231;
      8'b11101000 : _zz__zz_stateReg_75_34 = invSboxRom_232;
      8'b11101001 : _zz__zz_stateReg_75_34 = invSboxRom_233;
      8'b11101010 : _zz__zz_stateReg_75_34 = invSboxRom_234;
      8'b11101011 : _zz__zz_stateReg_75_34 = invSboxRom_235;
      8'b11101100 : _zz__zz_stateReg_75_34 = invSboxRom_236;
      8'b11101101 : _zz__zz_stateReg_75_34 = invSboxRom_237;
      8'b11101110 : _zz__zz_stateReg_75_34 = invSboxRom_238;
      8'b11101111 : _zz__zz_stateReg_75_34 = invSboxRom_239;
      8'b11110000 : _zz__zz_stateReg_75_34 = invSboxRom_240;
      8'b11110001 : _zz__zz_stateReg_75_34 = invSboxRom_241;
      8'b11110010 : _zz__zz_stateReg_75_34 = invSboxRom_242;
      8'b11110011 : _zz__zz_stateReg_75_34 = invSboxRom_243;
      8'b11110100 : _zz__zz_stateReg_75_34 = invSboxRom_244;
      8'b11110101 : _zz__zz_stateReg_75_34 = invSboxRom_245;
      8'b11110110 : _zz__zz_stateReg_75_34 = invSboxRom_246;
      8'b11110111 : _zz__zz_stateReg_75_34 = invSboxRom_247;
      8'b11111000 : _zz__zz_stateReg_75_34 = invSboxRom_248;
      8'b11111001 : _zz__zz_stateReg_75_34 = invSboxRom_249;
      8'b11111010 : _zz__zz_stateReg_75_34 = invSboxRom_250;
      8'b11111011 : _zz__zz_stateReg_75_34 = invSboxRom_251;
      8'b11111100 : _zz__zz_stateReg_75_34 = invSboxRom_252;
      8'b11111101 : _zz__zz_stateReg_75_34 = invSboxRom_253;
      8'b11111110 : _zz__zz_stateReg_75_34 = invSboxRom_254;
      default : _zz__zz_stateReg_75_34 = invSboxRom_255;
    endcase
  end

  assign rcon_0 = 8'h01;
  assign rcon_1 = 8'h02;
  assign rcon_2 = 8'h04;
  assign rcon_3 = 8'h08;
  assign rcon_4 = 8'h10;
  assign rcon_5 = 8'h20;
  assign rcon_6 = 8'h40;
  assign rcon_7 = 8'h80;
  assign rcon_8 = 8'h1b;
  assign rcon_9 = 8'h36;
  assign sboxRom_0 = 8'h63;
  assign sboxRom_1 = 8'h7c;
  assign sboxRom_2 = 8'h77;
  assign sboxRom_3 = 8'h7b;
  assign sboxRom_4 = 8'hf2;
  assign sboxRom_5 = 8'h6b;
  assign sboxRom_6 = 8'h6f;
  assign sboxRom_7 = 8'hc5;
  assign sboxRom_8 = 8'h30;
  assign sboxRom_9 = 8'h01;
  assign sboxRom_10 = 8'h67;
  assign sboxRom_11 = 8'h2b;
  assign sboxRom_12 = 8'hfe;
  assign sboxRom_13 = 8'hd7;
  assign sboxRom_14 = 8'hab;
  assign sboxRom_15 = 8'h76;
  assign sboxRom_16 = 8'hca;
  assign sboxRom_17 = 8'h82;
  assign sboxRom_18 = 8'hc9;
  assign sboxRom_19 = 8'h7d;
  assign sboxRom_20 = 8'hfa;
  assign sboxRom_21 = 8'h59;
  assign sboxRom_22 = 8'h47;
  assign sboxRom_23 = 8'hf0;
  assign sboxRom_24 = 8'had;
  assign sboxRom_25 = 8'hd4;
  assign sboxRom_26 = 8'ha2;
  assign sboxRom_27 = 8'haf;
  assign sboxRom_28 = 8'h9c;
  assign sboxRom_29 = 8'ha4;
  assign sboxRom_30 = 8'h72;
  assign sboxRom_31 = 8'hc0;
  assign sboxRom_32 = 8'hb7;
  assign sboxRom_33 = 8'hfd;
  assign sboxRom_34 = 8'h93;
  assign sboxRom_35 = 8'h26;
  assign sboxRom_36 = 8'h36;
  assign sboxRom_37 = 8'h3f;
  assign sboxRom_38 = 8'hf7;
  assign sboxRom_39 = 8'hcc;
  assign sboxRom_40 = 8'h34;
  assign sboxRom_41 = 8'ha5;
  assign sboxRom_42 = 8'he5;
  assign sboxRom_43 = 8'hf1;
  assign sboxRom_44 = 8'h71;
  assign sboxRom_45 = 8'hd8;
  assign sboxRom_46 = 8'h31;
  assign sboxRom_47 = 8'h15;
  assign sboxRom_48 = 8'h04;
  assign sboxRom_49 = 8'hc7;
  assign sboxRom_50 = 8'h23;
  assign sboxRom_51 = 8'hc3;
  assign sboxRom_52 = 8'h18;
  assign sboxRom_53 = 8'h96;
  assign sboxRom_54 = 8'h05;
  assign sboxRom_55 = 8'h9a;
  assign sboxRom_56 = 8'h07;
  assign sboxRom_57 = 8'h12;
  assign sboxRom_58 = 8'h80;
  assign sboxRom_59 = 8'he2;
  assign sboxRom_60 = 8'heb;
  assign sboxRom_61 = 8'h27;
  assign sboxRom_62 = 8'hb2;
  assign sboxRom_63 = 8'h75;
  assign sboxRom_64 = 8'h09;
  assign sboxRom_65 = 8'h83;
  assign sboxRom_66 = 8'h2c;
  assign sboxRom_67 = 8'h1a;
  assign sboxRom_68 = 8'h1b;
  assign sboxRom_69 = 8'h6e;
  assign sboxRom_70 = 8'h5a;
  assign sboxRom_71 = 8'ha0;
  assign sboxRom_72 = 8'h52;
  assign sboxRom_73 = 8'h3b;
  assign sboxRom_74 = 8'hd6;
  assign sboxRom_75 = 8'hb3;
  assign sboxRom_76 = 8'h29;
  assign sboxRom_77 = 8'he3;
  assign sboxRom_78 = 8'h2f;
  assign sboxRom_79 = 8'h84;
  assign sboxRom_80 = 8'h53;
  assign sboxRom_81 = 8'hd1;
  assign sboxRom_82 = 8'h0;
  assign sboxRom_83 = 8'hed;
  assign sboxRom_84 = 8'h20;
  assign sboxRom_85 = 8'hfc;
  assign sboxRom_86 = 8'hb1;
  assign sboxRom_87 = 8'h5b;
  assign sboxRom_88 = 8'h6a;
  assign sboxRom_89 = 8'hcb;
  assign sboxRom_90 = 8'hbe;
  assign sboxRom_91 = 8'h39;
  assign sboxRom_92 = 8'h4a;
  assign sboxRom_93 = 8'h4c;
  assign sboxRom_94 = 8'h58;
  assign sboxRom_95 = 8'hcf;
  assign sboxRom_96 = 8'hd0;
  assign sboxRom_97 = 8'hef;
  assign sboxRom_98 = 8'haa;
  assign sboxRom_99 = 8'hfb;
  assign sboxRom_100 = 8'h43;
  assign sboxRom_101 = 8'h4d;
  assign sboxRom_102 = 8'h33;
  assign sboxRom_103 = 8'h85;
  assign sboxRom_104 = 8'h45;
  assign sboxRom_105 = 8'hf9;
  assign sboxRom_106 = 8'h02;
  assign sboxRom_107 = 8'h7f;
  assign sboxRom_108 = 8'h50;
  assign sboxRom_109 = 8'h3c;
  assign sboxRom_110 = 8'h9f;
  assign sboxRom_111 = 8'ha8;
  assign sboxRom_112 = 8'h51;
  assign sboxRom_113 = 8'ha3;
  assign sboxRom_114 = 8'h40;
  assign sboxRom_115 = 8'h8f;
  assign sboxRom_116 = 8'h92;
  assign sboxRom_117 = 8'h9d;
  assign sboxRom_118 = 8'h38;
  assign sboxRom_119 = 8'hf5;
  assign sboxRom_120 = 8'hbc;
  assign sboxRom_121 = 8'hb6;
  assign sboxRom_122 = 8'hda;
  assign sboxRom_123 = 8'h21;
  assign sboxRom_124 = 8'h10;
  assign sboxRom_125 = 8'hff;
  assign sboxRom_126 = 8'hf3;
  assign sboxRom_127 = 8'hd2;
  assign sboxRom_128 = 8'hcd;
  assign sboxRom_129 = 8'h0c;
  assign sboxRom_130 = 8'h13;
  assign sboxRom_131 = 8'hec;
  assign sboxRom_132 = 8'h5f;
  assign sboxRom_133 = 8'h97;
  assign sboxRom_134 = 8'h44;
  assign sboxRom_135 = 8'h17;
  assign sboxRom_136 = 8'hc4;
  assign sboxRom_137 = 8'ha7;
  assign sboxRom_138 = 8'h7e;
  assign sboxRom_139 = 8'h3d;
  assign sboxRom_140 = 8'h64;
  assign sboxRom_141 = 8'h5d;
  assign sboxRom_142 = 8'h19;
  assign sboxRom_143 = 8'h73;
  assign sboxRom_144 = 8'h60;
  assign sboxRom_145 = 8'h81;
  assign sboxRom_146 = 8'h4f;
  assign sboxRom_147 = 8'hdc;
  assign sboxRom_148 = 8'h22;
  assign sboxRom_149 = 8'h2a;
  assign sboxRom_150 = 8'h90;
  assign sboxRom_151 = 8'h88;
  assign sboxRom_152 = 8'h46;
  assign sboxRom_153 = 8'hee;
  assign sboxRom_154 = 8'hb8;
  assign sboxRom_155 = 8'h14;
  assign sboxRom_156 = 8'hde;
  assign sboxRom_157 = 8'h5e;
  assign sboxRom_158 = 8'h0b;
  assign sboxRom_159 = 8'hdb;
  assign sboxRom_160 = 8'he0;
  assign sboxRom_161 = 8'h32;
  assign sboxRom_162 = 8'h3a;
  assign sboxRom_163 = 8'h0a;
  assign sboxRom_164 = 8'h49;
  assign sboxRom_165 = 8'h06;
  assign sboxRom_166 = 8'h24;
  assign sboxRom_167 = 8'h5c;
  assign sboxRom_168 = 8'hc2;
  assign sboxRom_169 = 8'hd3;
  assign sboxRom_170 = 8'hac;
  assign sboxRom_171 = 8'h62;
  assign sboxRom_172 = 8'h91;
  assign sboxRom_173 = 8'h95;
  assign sboxRom_174 = 8'he4;
  assign sboxRom_175 = 8'h79;
  assign sboxRom_176 = 8'he7;
  assign sboxRom_177 = 8'hc8;
  assign sboxRom_178 = 8'h37;
  assign sboxRom_179 = 8'h6d;
  assign sboxRom_180 = 8'h8d;
  assign sboxRom_181 = 8'hd5;
  assign sboxRom_182 = 8'h4e;
  assign sboxRom_183 = 8'ha9;
  assign sboxRom_184 = 8'h6c;
  assign sboxRom_185 = 8'h56;
  assign sboxRom_186 = 8'hf4;
  assign sboxRom_187 = 8'hea;
  assign sboxRom_188 = 8'h65;
  assign sboxRom_189 = 8'h7a;
  assign sboxRom_190 = 8'hae;
  assign sboxRom_191 = 8'h08;
  assign sboxRom_192 = 8'hba;
  assign sboxRom_193 = 8'h78;
  assign sboxRom_194 = 8'h25;
  assign sboxRom_195 = 8'h2e;
  assign sboxRom_196 = 8'h1c;
  assign sboxRom_197 = 8'ha6;
  assign sboxRom_198 = 8'hb4;
  assign sboxRom_199 = 8'hc6;
  assign sboxRom_200 = 8'he8;
  assign sboxRom_201 = 8'hdd;
  assign sboxRom_202 = 8'h74;
  assign sboxRom_203 = 8'h1f;
  assign sboxRom_204 = 8'h4b;
  assign sboxRom_205 = 8'hbd;
  assign sboxRom_206 = 8'h8b;
  assign sboxRom_207 = 8'h8a;
  assign sboxRom_208 = 8'h70;
  assign sboxRom_209 = 8'h3e;
  assign sboxRom_210 = 8'hb5;
  assign sboxRom_211 = 8'h66;
  assign sboxRom_212 = 8'h48;
  assign sboxRom_213 = 8'h03;
  assign sboxRom_214 = 8'hf6;
  assign sboxRom_215 = 8'h0e;
  assign sboxRom_216 = 8'h61;
  assign sboxRom_217 = 8'h35;
  assign sboxRom_218 = 8'h57;
  assign sboxRom_219 = 8'hb9;
  assign sboxRom_220 = 8'h86;
  assign sboxRom_221 = 8'hc1;
  assign sboxRom_222 = 8'h1d;
  assign sboxRom_223 = 8'h9e;
  assign sboxRom_224 = 8'he1;
  assign sboxRom_225 = 8'hf8;
  assign sboxRom_226 = 8'h98;
  assign sboxRom_227 = 8'h11;
  assign sboxRom_228 = 8'h69;
  assign sboxRom_229 = 8'hd9;
  assign sboxRom_230 = 8'h8e;
  assign sboxRom_231 = 8'h94;
  assign sboxRom_232 = 8'h9b;
  assign sboxRom_233 = 8'h1e;
  assign sboxRom_234 = 8'h87;
  assign sboxRom_235 = 8'he9;
  assign sboxRom_236 = 8'hce;
  assign sboxRom_237 = 8'h55;
  assign sboxRom_238 = 8'h28;
  assign sboxRom_239 = 8'hdf;
  assign sboxRom_240 = 8'h8c;
  assign sboxRom_241 = 8'ha1;
  assign sboxRom_242 = 8'h89;
  assign sboxRom_243 = 8'h0d;
  assign sboxRom_244 = 8'hbf;
  assign sboxRom_245 = 8'he6;
  assign sboxRom_246 = 8'h42;
  assign sboxRom_247 = 8'h68;
  assign sboxRom_248 = 8'h41;
  assign sboxRom_249 = 8'h99;
  assign sboxRom_250 = 8'h2d;
  assign sboxRom_251 = 8'h0f;
  assign sboxRom_252 = 8'hb0;
  assign sboxRom_253 = 8'h54;
  assign sboxRom_254 = 8'hbb;
  assign sboxRom_255 = 8'h16;
  assign invSboxRom_0 = 8'h52;
  assign invSboxRom_1 = 8'h09;
  assign invSboxRom_2 = 8'h6a;
  assign invSboxRom_3 = 8'hd5;
  assign invSboxRom_4 = 8'h30;
  assign invSboxRom_5 = 8'h36;
  assign invSboxRom_6 = 8'ha5;
  assign invSboxRom_7 = 8'h38;
  assign invSboxRom_8 = 8'hbf;
  assign invSboxRom_9 = 8'h40;
  assign invSboxRom_10 = 8'ha3;
  assign invSboxRom_11 = 8'h9e;
  assign invSboxRom_12 = 8'h81;
  assign invSboxRom_13 = 8'hf3;
  assign invSboxRom_14 = 8'hd7;
  assign invSboxRom_15 = 8'hfb;
  assign invSboxRom_16 = 8'h7c;
  assign invSboxRom_17 = 8'he3;
  assign invSboxRom_18 = 8'h39;
  assign invSboxRom_19 = 8'h82;
  assign invSboxRom_20 = 8'h9b;
  assign invSboxRom_21 = 8'h2f;
  assign invSboxRom_22 = 8'hff;
  assign invSboxRom_23 = 8'h87;
  assign invSboxRom_24 = 8'h34;
  assign invSboxRom_25 = 8'h8e;
  assign invSboxRom_26 = 8'h43;
  assign invSboxRom_27 = 8'h44;
  assign invSboxRom_28 = 8'hc4;
  assign invSboxRom_29 = 8'hde;
  assign invSboxRom_30 = 8'he9;
  assign invSboxRom_31 = 8'hcb;
  assign invSboxRom_32 = 8'h54;
  assign invSboxRom_33 = 8'h7b;
  assign invSboxRom_34 = 8'h94;
  assign invSboxRom_35 = 8'h32;
  assign invSboxRom_36 = 8'ha6;
  assign invSboxRom_37 = 8'hc2;
  assign invSboxRom_38 = 8'h23;
  assign invSboxRom_39 = 8'h3d;
  assign invSboxRom_40 = 8'hee;
  assign invSboxRom_41 = 8'h4c;
  assign invSboxRom_42 = 8'h95;
  assign invSboxRom_43 = 8'h0b;
  assign invSboxRom_44 = 8'h42;
  assign invSboxRom_45 = 8'hfa;
  assign invSboxRom_46 = 8'hc3;
  assign invSboxRom_47 = 8'h4e;
  assign invSboxRom_48 = 8'h08;
  assign invSboxRom_49 = 8'h2e;
  assign invSboxRom_50 = 8'ha1;
  assign invSboxRom_51 = 8'h66;
  assign invSboxRom_52 = 8'h28;
  assign invSboxRom_53 = 8'hd9;
  assign invSboxRom_54 = 8'h24;
  assign invSboxRom_55 = 8'hb2;
  assign invSboxRom_56 = 8'h76;
  assign invSboxRom_57 = 8'h5b;
  assign invSboxRom_58 = 8'ha2;
  assign invSboxRom_59 = 8'h49;
  assign invSboxRom_60 = 8'h6d;
  assign invSboxRom_61 = 8'h8b;
  assign invSboxRom_62 = 8'hd1;
  assign invSboxRom_63 = 8'h25;
  assign invSboxRom_64 = 8'h72;
  assign invSboxRom_65 = 8'hf8;
  assign invSboxRom_66 = 8'hf6;
  assign invSboxRom_67 = 8'h64;
  assign invSboxRom_68 = 8'h86;
  assign invSboxRom_69 = 8'h68;
  assign invSboxRom_70 = 8'h98;
  assign invSboxRom_71 = 8'h16;
  assign invSboxRom_72 = 8'hd4;
  assign invSboxRom_73 = 8'ha4;
  assign invSboxRom_74 = 8'h5c;
  assign invSboxRom_75 = 8'hcc;
  assign invSboxRom_76 = 8'h5d;
  assign invSboxRom_77 = 8'h65;
  assign invSboxRom_78 = 8'hb6;
  assign invSboxRom_79 = 8'h92;
  assign invSboxRom_80 = 8'h6c;
  assign invSboxRom_81 = 8'h70;
  assign invSboxRom_82 = 8'h48;
  assign invSboxRom_83 = 8'h50;
  assign invSboxRom_84 = 8'hfd;
  assign invSboxRom_85 = 8'hed;
  assign invSboxRom_86 = 8'hb9;
  assign invSboxRom_87 = 8'hda;
  assign invSboxRom_88 = 8'h5e;
  assign invSboxRom_89 = 8'h15;
  assign invSboxRom_90 = 8'h46;
  assign invSboxRom_91 = 8'h57;
  assign invSboxRom_92 = 8'ha7;
  assign invSboxRom_93 = 8'h8d;
  assign invSboxRom_94 = 8'h9d;
  assign invSboxRom_95 = 8'h84;
  assign invSboxRom_96 = 8'h90;
  assign invSboxRom_97 = 8'hd8;
  assign invSboxRom_98 = 8'hab;
  assign invSboxRom_99 = 8'h0;
  assign invSboxRom_100 = 8'h8c;
  assign invSboxRom_101 = 8'hbc;
  assign invSboxRom_102 = 8'hd3;
  assign invSboxRom_103 = 8'h0a;
  assign invSboxRom_104 = 8'hf7;
  assign invSboxRom_105 = 8'he4;
  assign invSboxRom_106 = 8'h58;
  assign invSboxRom_107 = 8'h05;
  assign invSboxRom_108 = 8'hb8;
  assign invSboxRom_109 = 8'hb3;
  assign invSboxRom_110 = 8'h45;
  assign invSboxRom_111 = 8'h06;
  assign invSboxRom_112 = 8'hd0;
  assign invSboxRom_113 = 8'h2c;
  assign invSboxRom_114 = 8'h1e;
  assign invSboxRom_115 = 8'h8f;
  assign invSboxRom_116 = 8'hca;
  assign invSboxRom_117 = 8'h3f;
  assign invSboxRom_118 = 8'h0f;
  assign invSboxRom_119 = 8'h02;
  assign invSboxRom_120 = 8'hc1;
  assign invSboxRom_121 = 8'haf;
  assign invSboxRom_122 = 8'hbd;
  assign invSboxRom_123 = 8'h03;
  assign invSboxRom_124 = 8'h01;
  assign invSboxRom_125 = 8'h13;
  assign invSboxRom_126 = 8'h8a;
  assign invSboxRom_127 = 8'h6b;
  assign invSboxRom_128 = 8'h3a;
  assign invSboxRom_129 = 8'h91;
  assign invSboxRom_130 = 8'h11;
  assign invSboxRom_131 = 8'h41;
  assign invSboxRom_132 = 8'h4f;
  assign invSboxRom_133 = 8'h67;
  assign invSboxRom_134 = 8'hdc;
  assign invSboxRom_135 = 8'hea;
  assign invSboxRom_136 = 8'h97;
  assign invSboxRom_137 = 8'hf2;
  assign invSboxRom_138 = 8'hcf;
  assign invSboxRom_139 = 8'hce;
  assign invSboxRom_140 = 8'hf0;
  assign invSboxRom_141 = 8'hb4;
  assign invSboxRom_142 = 8'he6;
  assign invSboxRom_143 = 8'h73;
  assign invSboxRom_144 = 8'h96;
  assign invSboxRom_145 = 8'hac;
  assign invSboxRom_146 = 8'h74;
  assign invSboxRom_147 = 8'h22;
  assign invSboxRom_148 = 8'he7;
  assign invSboxRom_149 = 8'had;
  assign invSboxRom_150 = 8'h35;
  assign invSboxRom_151 = 8'h85;
  assign invSboxRom_152 = 8'he2;
  assign invSboxRom_153 = 8'hf9;
  assign invSboxRom_154 = 8'h37;
  assign invSboxRom_155 = 8'he8;
  assign invSboxRom_156 = 8'h1c;
  assign invSboxRom_157 = 8'h75;
  assign invSboxRom_158 = 8'hdf;
  assign invSboxRom_159 = 8'h6e;
  assign invSboxRom_160 = 8'h47;
  assign invSboxRom_161 = 8'hf1;
  assign invSboxRom_162 = 8'h1a;
  assign invSboxRom_163 = 8'h71;
  assign invSboxRom_164 = 8'h1d;
  assign invSboxRom_165 = 8'h29;
  assign invSboxRom_166 = 8'hc5;
  assign invSboxRom_167 = 8'h89;
  assign invSboxRom_168 = 8'h6f;
  assign invSboxRom_169 = 8'hb7;
  assign invSboxRom_170 = 8'h62;
  assign invSboxRom_171 = 8'h0e;
  assign invSboxRom_172 = 8'haa;
  assign invSboxRom_173 = 8'h18;
  assign invSboxRom_174 = 8'hbe;
  assign invSboxRom_175 = 8'h1b;
  assign invSboxRom_176 = 8'hfc;
  assign invSboxRom_177 = 8'h56;
  assign invSboxRom_178 = 8'h3e;
  assign invSboxRom_179 = 8'h4b;
  assign invSboxRom_180 = 8'hc6;
  assign invSboxRom_181 = 8'hd2;
  assign invSboxRom_182 = 8'h79;
  assign invSboxRom_183 = 8'h20;
  assign invSboxRom_184 = 8'h9a;
  assign invSboxRom_185 = 8'hdb;
  assign invSboxRom_186 = 8'hc0;
  assign invSboxRom_187 = 8'hfe;
  assign invSboxRom_188 = 8'h78;
  assign invSboxRom_189 = 8'hcd;
  assign invSboxRom_190 = 8'h5a;
  assign invSboxRom_191 = 8'hf4;
  assign invSboxRom_192 = 8'h1f;
  assign invSboxRom_193 = 8'hdd;
  assign invSboxRom_194 = 8'ha8;
  assign invSboxRom_195 = 8'h33;
  assign invSboxRom_196 = 8'h88;
  assign invSboxRom_197 = 8'h07;
  assign invSboxRom_198 = 8'hc7;
  assign invSboxRom_199 = 8'h31;
  assign invSboxRom_200 = 8'hb1;
  assign invSboxRom_201 = 8'h12;
  assign invSboxRom_202 = 8'h10;
  assign invSboxRom_203 = 8'h59;
  assign invSboxRom_204 = 8'h27;
  assign invSboxRom_205 = 8'h80;
  assign invSboxRom_206 = 8'hec;
  assign invSboxRom_207 = 8'h5f;
  assign invSboxRom_208 = 8'h60;
  assign invSboxRom_209 = 8'h51;
  assign invSboxRom_210 = 8'h7f;
  assign invSboxRom_211 = 8'ha9;
  assign invSboxRom_212 = 8'h19;
  assign invSboxRom_213 = 8'hb5;
  assign invSboxRom_214 = 8'h4a;
  assign invSboxRom_215 = 8'h0d;
  assign invSboxRom_216 = 8'h2d;
  assign invSboxRom_217 = 8'he5;
  assign invSboxRom_218 = 8'h7a;
  assign invSboxRom_219 = 8'h9f;
  assign invSboxRom_220 = 8'h93;
  assign invSboxRom_221 = 8'hc9;
  assign invSboxRom_222 = 8'h9c;
  assign invSboxRom_223 = 8'hef;
  assign invSboxRom_224 = 8'ha0;
  assign invSboxRom_225 = 8'he0;
  assign invSboxRom_226 = 8'h3b;
  assign invSboxRom_227 = 8'h4d;
  assign invSboxRom_228 = 8'hae;
  assign invSboxRom_229 = 8'h2a;
  assign invSboxRom_230 = 8'hf5;
  assign invSboxRom_231 = 8'hb0;
  assign invSboxRom_232 = 8'hc8;
  assign invSboxRom_233 = 8'heb;
  assign invSboxRom_234 = 8'hbb;
  assign invSboxRom_235 = 8'h3c;
  assign invSboxRom_236 = 8'h83;
  assign invSboxRom_237 = 8'h53;
  assign invSboxRom_238 = 8'h99;
  assign invSboxRom_239 = 8'h61;
  assign invSboxRom_240 = 8'h17;
  assign invSboxRom_241 = 8'h2b;
  assign invSboxRom_242 = 8'h04;
  assign invSboxRom_243 = 8'h7e;
  assign invSboxRom_244 = 8'hba;
  assign invSboxRom_245 = 8'h77;
  assign invSboxRom_246 = 8'hd6;
  assign invSboxRom_247 = 8'h26;
  assign invSboxRom_248 = 8'he1;
  assign invSboxRom_249 = 8'h69;
  assign invSboxRom_250 = 8'h14;
  assign invSboxRom_251 = 8'h63;
  assign invSboxRom_252 = 8'h55;
  assign invSboxRom_253 = 8'h21;
  assign invSboxRom_254 = 8'h0c;
  assign invSboxRom_255 = 8'h7d;
  assign io_busy = running;
  always @(*) begin
    io_done = 1'b0;
    if(!when_AES128_l215) begin
      if(when_AES128_l229) begin
        if(when_AES128_l291) begin
          io_done = 1'b1;
        end
      end else begin
        if(!when_AES128_l299) begin
          if(!precomputeRunning) begin
            if(when_AES128_l324) begin
              if(when_AES128_l383) begin
                io_done = 1'b1;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    io_dataOut = stateReg;
    if(!when_AES128_l215) begin
      if(when_AES128_l229) begin
        if(when_AES128_l291) begin
          io_dataOut = stateReg;
        end
      end else begin
        if(!when_AES128_l299) begin
          if(!precomputeRunning) begin
            if(when_AES128_l324) begin
              if(when_AES128_l383) begin
                io_dataOut = stateReg;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    newStateComb = 128'h0;
    if(!when_AES128_l215) begin
      if(when_AES128_l229) begin
        newStateComb = _zz_stateReg_68;
      end
    end
  end

  always @(*) begin
    rkBitsUsedComb = 128'h0;
    if(!when_AES128_l215) begin
      if(when_AES128_l229) begin
        rkBitsUsedComb = _zz_stateReg_69;
      end
    end
  end

  assign when_AES128_l215 = ((io_start && (! running)) && (! io_decrypt));
  assign _zz_stateReg = io_key[127 : 96];
  assign _zz_stateReg_1 = io_key[95 : 64];
  assign _zz_stateReg_2 = io_key[63 : 32];
  assign _zz_stateReg_3 = io_key[31 : 0];
  assign _zz_stateReg_4 = _zz__zz_stateReg_4;
  assign _zz_stateReg_8 = _zz__zz_stateReg_8;
  assign _zz_stateReg_12 = _zz__zz_stateReg_12;
  assign _zz_stateReg_16 = _zz__zz_stateReg_16;
  assign _zz_stateReg_5 = _zz__zz_stateReg_5;
  assign _zz_stateReg_9 = _zz__zz_stateReg_9;
  assign _zz_stateReg_13 = _zz__zz_stateReg_13;
  assign _zz_stateReg_17 = _zz__zz_stateReg_17;
  assign _zz_stateReg_6 = _zz__zz_stateReg_6;
  assign _zz_stateReg_10 = _zz__zz_stateReg_10;
  assign _zz_stateReg_14 = _zz__zz_stateReg_14;
  assign _zz_stateReg_18 = _zz__zz_stateReg_18;
  assign _zz_stateReg_7 = _zz__zz_stateReg_7;
  assign _zz_stateReg_11 = _zz__zz_stateReg_11;
  assign _zz_stateReg_15 = _zz__zz_stateReg_15;
  assign _zz_stateReg_19 = _zz__zz_stateReg_19;
  assign when_AES128_l257 = (roundCount == 4'b1001);
  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_20 = _zz_stateReg_4;
    end else begin
      _zz_stateReg_20 = ((((_zz_stateReg_4[7] ? (_zz_stateReg_36 ^ 8'h1b) : _zz_stateReg_36) ^ ((_zz_stateReg_5[7] ? (_zz_stateReg_37 ^ 8'h1b) : _zz_stateReg_37) ^ _zz_stateReg_5)) ^ _zz_stateReg_6) ^ _zz_stateReg_7);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_21 = _zz_stateReg_5;
    end else begin
      _zz_stateReg_21 = (((_zz_stateReg_4 ^ (_zz_stateReg_5[7] ? (_zz_stateReg_38 ^ 8'h1b) : _zz_stateReg_38)) ^ ((_zz_stateReg_6[7] ? (_zz_stateReg_39 ^ 8'h1b) : _zz_stateReg_39) ^ _zz_stateReg_6)) ^ _zz_stateReg_7);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_22 = _zz_stateReg_6;
    end else begin
      _zz_stateReg_22 = (((_zz_stateReg_4 ^ _zz_stateReg_5) ^ (_zz_stateReg_6[7] ? (_zz_stateReg_40 ^ 8'h1b) : _zz_stateReg_40)) ^ ((_zz_stateReg_7[7] ? (_zz_stateReg_41 ^ 8'h1b) : _zz_stateReg_41) ^ _zz_stateReg_7));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_23 = _zz_stateReg_7;
    end else begin
      _zz_stateReg_23 = (((((_zz_stateReg_4[7] ? (_zz_stateReg_42 ^ 8'h1b) : _zz_stateReg_42) ^ _zz_stateReg_4) ^ _zz_stateReg_5) ^ _zz_stateReg_6) ^ (_zz_stateReg_7[7] ? (_zz_stateReg_43 ^ 8'h1b) : _zz_stateReg_43));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_24 = _zz_stateReg_8;
    end else begin
      _zz_stateReg_24 = ((((_zz_stateReg_8[7] ? (_zz_stateReg_44 ^ 8'h1b) : _zz_stateReg_44) ^ ((_zz_stateReg_9[7] ? (_zz_stateReg_45 ^ 8'h1b) : _zz_stateReg_45) ^ _zz_stateReg_9)) ^ _zz_stateReg_10) ^ _zz_stateReg_11);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_25 = _zz_stateReg_9;
    end else begin
      _zz_stateReg_25 = (((_zz_stateReg_8 ^ (_zz_stateReg_9[7] ? (_zz_stateReg_46 ^ 8'h1b) : _zz_stateReg_46)) ^ ((_zz_stateReg_10[7] ? (_zz_stateReg_47 ^ 8'h1b) : _zz_stateReg_47) ^ _zz_stateReg_10)) ^ _zz_stateReg_11);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_26 = _zz_stateReg_10;
    end else begin
      _zz_stateReg_26 = (((_zz_stateReg_8 ^ _zz_stateReg_9) ^ (_zz_stateReg_10[7] ? (_zz_stateReg_48 ^ 8'h1b) : _zz_stateReg_48)) ^ ((_zz_stateReg_11[7] ? (_zz_stateReg_49 ^ 8'h1b) : _zz_stateReg_49) ^ _zz_stateReg_11));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_27 = _zz_stateReg_11;
    end else begin
      _zz_stateReg_27 = (((((_zz_stateReg_8[7] ? (_zz_stateReg_50 ^ 8'h1b) : _zz_stateReg_50) ^ _zz_stateReg_8) ^ _zz_stateReg_9) ^ _zz_stateReg_10) ^ (_zz_stateReg_11[7] ? (_zz_stateReg_51 ^ 8'h1b) : _zz_stateReg_51));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_28 = _zz_stateReg_12;
    end else begin
      _zz_stateReg_28 = ((((_zz_stateReg_12[7] ? (_zz_stateReg_52 ^ 8'h1b) : _zz_stateReg_52) ^ ((_zz_stateReg_13[7] ? (_zz_stateReg_53 ^ 8'h1b) : _zz_stateReg_53) ^ _zz_stateReg_13)) ^ _zz_stateReg_14) ^ _zz_stateReg_15);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_29 = _zz_stateReg_13;
    end else begin
      _zz_stateReg_29 = (((_zz_stateReg_12 ^ (_zz_stateReg_13[7] ? (_zz_stateReg_54 ^ 8'h1b) : _zz_stateReg_54)) ^ ((_zz_stateReg_14[7] ? (_zz_stateReg_55 ^ 8'h1b) : _zz_stateReg_55) ^ _zz_stateReg_14)) ^ _zz_stateReg_15);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_30 = _zz_stateReg_14;
    end else begin
      _zz_stateReg_30 = (((_zz_stateReg_12 ^ _zz_stateReg_13) ^ (_zz_stateReg_14[7] ? (_zz_stateReg_56 ^ 8'h1b) : _zz_stateReg_56)) ^ ((_zz_stateReg_15[7] ? (_zz_stateReg_57 ^ 8'h1b) : _zz_stateReg_57) ^ _zz_stateReg_15));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_31 = _zz_stateReg_15;
    end else begin
      _zz_stateReg_31 = (((((_zz_stateReg_12[7] ? (_zz_stateReg_58 ^ 8'h1b) : _zz_stateReg_58) ^ _zz_stateReg_12) ^ _zz_stateReg_13) ^ _zz_stateReg_14) ^ (_zz_stateReg_15[7] ? (_zz_stateReg_59 ^ 8'h1b) : _zz_stateReg_59));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_32 = _zz_stateReg_16;
    end else begin
      _zz_stateReg_32 = ((((_zz_stateReg_16[7] ? (_zz_stateReg_60 ^ 8'h1b) : _zz_stateReg_60) ^ ((_zz_stateReg_17[7] ? (_zz_stateReg_61 ^ 8'h1b) : _zz_stateReg_61) ^ _zz_stateReg_17)) ^ _zz_stateReg_18) ^ _zz_stateReg_19);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_33 = _zz_stateReg_17;
    end else begin
      _zz_stateReg_33 = (((_zz_stateReg_16 ^ (_zz_stateReg_17[7] ? (_zz_stateReg_62 ^ 8'h1b) : _zz_stateReg_62)) ^ ((_zz_stateReg_18[7] ? (_zz_stateReg_63 ^ 8'h1b) : _zz_stateReg_63) ^ _zz_stateReg_18)) ^ _zz_stateReg_19);
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_34 = _zz_stateReg_18;
    end else begin
      _zz_stateReg_34 = (((_zz_stateReg_16 ^ _zz_stateReg_17) ^ (_zz_stateReg_18[7] ? (_zz_stateReg_64 ^ 8'h1b) : _zz_stateReg_64)) ^ ((_zz_stateReg_19[7] ? (_zz_stateReg_65 ^ 8'h1b) : _zz_stateReg_65) ^ _zz_stateReg_19));
    end
  end

  always @(*) begin
    if(when_AES128_l257) begin
      _zz_stateReg_35 = _zz_stateReg_19;
    end else begin
      _zz_stateReg_35 = (((((_zz_stateReg_16[7] ? (_zz_stateReg_66 ^ 8'h1b) : _zz_stateReg_66) ^ _zz_stateReg_16) ^ _zz_stateReg_17) ^ _zz_stateReg_18) ^ (_zz_stateReg_19[7] ? (_zz_stateReg_67 ^ 8'h1b) : _zz_stateReg_67));
    end
  end

  assign _zz_stateReg_36 = _zz__zz_stateReg_36[7 : 0];
  assign _zz_stateReg_37 = _zz__zz_stateReg_37[7 : 0];
  assign _zz_stateReg_38 = _zz__zz_stateReg_38[7 : 0];
  assign _zz_stateReg_39 = _zz__zz_stateReg_39[7 : 0];
  assign _zz_stateReg_40 = _zz__zz_stateReg_40[7 : 0];
  assign _zz_stateReg_41 = _zz__zz_stateReg_41[7 : 0];
  assign _zz_stateReg_42 = _zz__zz_stateReg_42[7 : 0];
  assign _zz_stateReg_43 = _zz__zz_stateReg_43[7 : 0];
  assign _zz_stateReg_44 = _zz__zz_stateReg_44[7 : 0];
  assign _zz_stateReg_45 = _zz__zz_stateReg_45[7 : 0];
  assign _zz_stateReg_46 = _zz__zz_stateReg_46[7 : 0];
  assign _zz_stateReg_47 = _zz__zz_stateReg_47[7 : 0];
  assign _zz_stateReg_48 = _zz__zz_stateReg_48[7 : 0];
  assign _zz_stateReg_49 = _zz__zz_stateReg_49[7 : 0];
  assign _zz_stateReg_50 = _zz__zz_stateReg_50[7 : 0];
  assign _zz_stateReg_51 = _zz__zz_stateReg_51[7 : 0];
  assign _zz_stateReg_52 = _zz__zz_stateReg_52[7 : 0];
  assign _zz_stateReg_53 = _zz__zz_stateReg_53[7 : 0];
  assign _zz_stateReg_54 = _zz__zz_stateReg_54[7 : 0];
  assign _zz_stateReg_55 = _zz__zz_stateReg_55[7 : 0];
  assign _zz_stateReg_56 = _zz__zz_stateReg_56[7 : 0];
  assign _zz_stateReg_57 = _zz__zz_stateReg_57[7 : 0];
  assign _zz_stateReg_58 = _zz__zz_stateReg_58[7 : 0];
  assign _zz_stateReg_59 = _zz__zz_stateReg_59[7 : 0];
  assign _zz_stateReg_60 = _zz__zz_stateReg_60[7 : 0];
  assign _zz_stateReg_61 = _zz__zz_stateReg_61[7 : 0];
  assign _zz_stateReg_62 = _zz__zz_stateReg_62[7 : 0];
  assign _zz_stateReg_63 = _zz__zz_stateReg_63[7 : 0];
  assign _zz_stateReg_64 = _zz__zz_stateReg_64[7 : 0];
  assign _zz_stateReg_65 = _zz__zz_stateReg_65[7 : 0];
  assign _zz_stateReg_66 = _zz__zz_stateReg_66[7 : 0];
  assign _zz_stateReg_67 = _zz__zz_stateReg_67[7 : 0];
  assign _zz_stateReg_68 = {{{{{{{{{{{_zz__zz_stateReg_68,_zz__zz_stateReg_68_1},_zz_stateReg_26},_zz_stateReg_27},_zz_stateReg_28},_zz_stateReg_29},_zz_stateReg_30},_zz_stateReg_31},_zz_stateReg_32},_zz_stateReg_33},_zz_stateReg_34},_zz_stateReg_35};
  assign _zz_roundKeyReg_0 = _zz__zz_roundKeyReg_0;
  assign _zz_roundKeyReg_0_1 = {roundKeyReg_3[23 : 0],roundKeyReg_3[31 : 24]};
  assign _zz_roundKeyReg_0_2 = (roundKeyReg_0 ^ ({{{_zz__zz_roundKeyReg_0_2,_zz__zz_roundKeyReg_0_2_2},_zz__zz_roundKeyReg_0_2_4},_zz__zz_roundKeyReg_0_2_6} ^ {_zz_roundKeyReg_0,24'h0}));
  assign _zz_roundKeyReg_1 = (roundKeyReg_1 ^ _zz_roundKeyReg_0_2);
  assign _zz_roundKeyReg_2 = (roundKeyReg_2 ^ _zz_roundKeyReg_1);
  assign _zz_roundKeyReg_3 = (roundKeyReg_3 ^ _zz_roundKeyReg_2);
  assign _zz_stateReg_69 = {{{{{{{{{_zz__zz_stateReg_69,_zz__zz_stateReg_69_1},_zz__zz_stateReg_69_2},_zz_roundKeyReg_2[23 : 16]},_zz_roundKeyReg_2[15 : 8]},_zz_roundKeyReg_2[7 : 0]},_zz_roundKeyReg_3[31 : 24]},_zz_roundKeyReg_3[23 : 16]},_zz_roundKeyReg_3[15 : 8]},_zz_roundKeyReg_3[7 : 0]};
  assign when_AES128_l291 = (roundCount == 4'b1010);
  assign when_AES128_l297 = (rconCounter < 4'b1001);
  assign _zz_stateReg_70 = {roundKeyReg_3[23 : 0],roundKeyReg_3[31 : 24]};
  assign _zz_stateReg_71 = (roundKeyReg_0 ^ ({{{_zz__zz_stateReg_71,_zz__zz_stateReg_71_2},_zz__zz_stateReg_71_4},_zz__zz_stateReg_71_6} ^ {_zz__zz_stateReg_71_8,24'h0}));
  assign _zz_stateReg_72 = (roundKeyReg_1 ^ _zz_stateReg_71);
  assign _zz_stateReg_73 = (roundKeyReg_2 ^ _zz_stateReg_72);
  assign _zz_stateReg_74 = (roundKeyReg_3 ^ _zz_stateReg_73);
  assign when_AES128_l313 = (precomputeCounter == 4'b1001);
  assign _zz_roundKeyReg_3_1 = (roundKeyReg_3 ^ roundKeyReg_2);
  assign _zz_roundKeyReg_2_1 = (roundKeyReg_2 ^ roundKeyReg_1);
  assign _zz_roundKeyReg_1_1 = (roundKeyReg_1 ^ roundKeyReg_0);
  assign _zz_roundKeyReg_0_3 = {_zz_roundKeyReg_3_1[23 : 0],_zz_roundKeyReg_3_1[31 : 24]};
  assign _zz_roundKeyReg_0_4 = (roundKeyReg_0 ^ ({{{_zz__zz_roundKeyReg_0_4,_zz__zz_roundKeyReg_0_4_2},_zz__zz_roundKeyReg_0_4_4},_zz__zz_roundKeyReg_0_4_6} ^ {_zz_roundKeyReg_0,24'h0}));
  assign _zz_stateReg_75 = ({{{{{{_zz__zz_stateReg_75,_zz__zz_stateReg_75_23},_zz__zz_stateReg_75_26},_zz__zz_stateReg_75_28},_zz__zz_stateReg_75_30},_zz__zz_stateReg_75_32},_zz__zz_stateReg_75_34} ^ {{{{{{_zz__zz_stateReg_75_36,_zz__zz_stateReg_75_40},_zz__zz_stateReg_75_41},_zz_roundKeyReg_3_1[31 : 24]},_zz_roundKeyReg_3_1[23 : 16]},_zz_roundKeyReg_3_1[15 : 8]},_zz_roundKeyReg_3_1[7 : 0]});
  assign _zz_stateReg_76 = _zz_stateReg_75[127 : 120];
  assign _zz_stateReg_77 = _zz_stateReg_75[119 : 112];
  assign _zz_stateReg_78 = _zz_stateReg_75[111 : 104];
  assign _zz_stateReg_79 = _zz_stateReg_75[103 : 96];
  assign _zz_stateReg_80 = _zz_stateReg_75[95 : 88];
  assign _zz_stateReg_81 = _zz_stateReg_75[87 : 80];
  assign _zz_stateReg_82 = _zz_stateReg_75[79 : 72];
  assign _zz_stateReg_83 = _zz_stateReg_75[71 : 64];
  assign _zz_stateReg_84 = _zz_stateReg_75[63 : 56];
  assign _zz_stateReg_85 = _zz_stateReg_75[55 : 48];
  assign _zz_stateReg_86 = _zz_stateReg_75[47 : 40];
  assign _zz_stateReg_87 = _zz_stateReg_75[39 : 32];
  assign _zz_stateReg_88 = _zz_stateReg_75[31 : 24];
  assign _zz_stateReg_89 = _zz_stateReg_75[23 : 16];
  assign _zz_stateReg_90 = _zz_stateReg_75[15 : 8];
  assign _zz_stateReg_91 = _zz_stateReg_75[7 : 0];
  always @(*) begin
    _zz_stateReg_92 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_92 = _zz_stateReg_76;
    end else begin
      _zz_stateReg_92 = (((((_zz__zz_stateReg_92 ^ _zz__zz_stateReg_92_1) ^ (_zz__zz_stateReg_92_2 ? _zz__zz_stateReg_92_3 : _zz_stateReg_116)) ^ ((_zz__zz_stateReg_92_4 ^ _zz__zz_stateReg_92_5) ^ _zz_stateReg_77)) ^ (((_zz__zz_stateReg_92_6 ? _zz__zz_stateReg_92_7 : _zz_stateReg_127) ^ (_zz__zz_stateReg_92_8 ? _zz__zz_stateReg_92_9 : _zz_stateReg_130)) ^ _zz_stateReg_78)) ^ ((_zz_stateReg_134[7] ? (_zz_stateReg_135 ^ 8'h1b) : _zz_stateReg_135) ^ _zz_stateReg_79));
    end
  end

  always @(*) begin
    _zz_stateReg_93 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_93 = _zz_stateReg_77;
    end else begin
      _zz_stateReg_93 = (((((_zz__zz_stateReg_93 ? _zz__zz_stateReg_93_1 : _zz_stateReg_140) ^ _zz_stateReg_76) ^ ((_zz__zz_stateReg_93_2 ^ _zz__zz_stateReg_93_3) ^ (_zz__zz_stateReg_93_4 ? _zz__zz_stateReg_93_5 : _zz_stateReg_149))) ^ (((_zz__zz_stateReg_93_6 ? _zz__zz_stateReg_93_7 : _zz_stateReg_154) ^ (_zz__zz_stateReg_93_8 ? _zz__zz_stateReg_93_9 : _zz_stateReg_155)) ^ _zz_stateReg_78)) ^ (((_zz_stateReg_159[7] ? (_zz_stateReg_160 ^ _zz__zz_stateReg_93_10) : _zz_stateReg_160) ^ (_zz_stateReg_162[7] ? (_zz_stateReg_163 ^ _zz__zz_stateReg_93_11) : _zz_stateReg_163)) ^ _zz_stateReg_79));
    end
  end

  always @(*) begin
    _zz_stateReg_94 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_94 = _zz_stateReg_78;
    end else begin
      _zz_stateReg_94 = (((((_zz__zz_stateReg_94 ^ _zz__zz_stateReg_94_1) ^ _zz_stateReg_76) ^ ((_zz__zz_stateReg_94_2 ? _zz__zz_stateReg_94_3 : _zz_stateReg_176) ^ _zz_stateReg_77)) ^ (((_zz__zz_stateReg_94_4 ? _zz__zz_stateReg_94_5 : _zz_stateReg_181) ^ (_zz__zz_stateReg_94_6 ? _zz__zz_stateReg_94_7 : _zz_stateReg_184)) ^ (_zz_stateReg_78[7] ? (_zz_stateReg_185 ^ _zz__zz_stateReg_94_8) : _zz_stateReg_185))) ^ (((_zz_stateReg_189[7] ? (_zz_stateReg_190 ^ _zz__zz_stateReg_94_9) : _zz_stateReg_190) ^ (_zz_stateReg_79[7] ? (_zz_stateReg_191 ^ _zz__zz_stateReg_94_10) : _zz_stateReg_191)) ^ _zz_stateReg_79));
    end
  end

  always @(*) begin
    _zz_stateReg_95 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_95 = _zz_stateReg_79;
    end else begin
      _zz_stateReg_95 = (((((_zz__zz_stateReg_95 ^ _zz__zz_stateReg_95_1) ^ _zz_stateReg_76) ^ ((_zz__zz_stateReg_95_2 ^ _zz__zz_stateReg_95_3) ^ _zz_stateReg_77)) ^ ((_zz_stateReg_209[7] ? (_zz_stateReg_210 ^ _zz__zz_stateReg_95_4) : _zz_stateReg_210) ^ _zz_stateReg_78)) ^ (((_zz_stateReg_214[7] ? (_zz_stateReg_215 ^ _zz__zz_stateReg_95_5) : _zz_stateReg_215) ^ (_zz_stateReg_217[7] ? (_zz_stateReg_218 ^ _zz__zz_stateReg_95_6) : _zz_stateReg_218)) ^ (_zz_stateReg_79[7] ? (_zz_stateReg_219 ^ 8'h1b) : _zz_stateReg_219)));
    end
  end

  always @(*) begin
    _zz_stateReg_96 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_96 = _zz_stateReg_80;
    end else begin
      _zz_stateReg_96 = (((((_zz__zz_stateReg_96 ^ _zz__zz_stateReg_96_1) ^ (_zz__zz_stateReg_96_2 ? _zz__zz_stateReg_96_3 : _zz_stateReg_228)) ^ ((_zz__zz_stateReg_96_4 ^ _zz__zz_stateReg_96_5) ^ _zz_stateReg_81)) ^ (((_zz__zz_stateReg_96_6 ? _zz__zz_stateReg_96_7 : _zz_stateReg_239) ^ (_zz__zz_stateReg_96_8 ? _zz__zz_stateReg_96_9 : _zz_stateReg_242)) ^ _zz_stateReg_82)) ^ ((_zz_stateReg_246[7] ? (_zz_stateReg_247 ^ 8'h1b) : _zz_stateReg_247) ^ _zz_stateReg_83));
    end
  end

  always @(*) begin
    _zz_stateReg_97 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_97 = _zz_stateReg_81;
    end else begin
      _zz_stateReg_97 = (((((_zz__zz_stateReg_97 ? _zz__zz_stateReg_97_1 : _zz_stateReg_252) ^ _zz_stateReg_80) ^ ((_zz__zz_stateReg_97_2 ^ _zz__zz_stateReg_97_3) ^ (_zz__zz_stateReg_97_4 ? _zz__zz_stateReg_97_5 : _zz_stateReg_261))) ^ (((_zz__zz_stateReg_97_6 ? _zz__zz_stateReg_97_7 : _zz_stateReg_266) ^ (_zz__zz_stateReg_97_8 ? _zz__zz_stateReg_97_9 : _zz_stateReg_267)) ^ _zz_stateReg_82)) ^ (((_zz_stateReg_271[7] ? (_zz_stateReg_272 ^ _zz__zz_stateReg_97_10) : _zz_stateReg_272) ^ (_zz_stateReg_274[7] ? (_zz_stateReg_275 ^ _zz__zz_stateReg_97_11) : _zz_stateReg_275)) ^ _zz_stateReg_83));
    end
  end

  always @(*) begin
    _zz_stateReg_98 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_98 = _zz_stateReg_82;
    end else begin
      _zz_stateReg_98 = (((((_zz__zz_stateReg_98 ^ _zz__zz_stateReg_98_1) ^ _zz_stateReg_80) ^ ((_zz__zz_stateReg_98_2 ? _zz__zz_stateReg_98_3 : _zz_stateReg_288) ^ _zz_stateReg_81)) ^ (((_zz__zz_stateReg_98_4 ? _zz__zz_stateReg_98_5 : _zz_stateReg_293) ^ (_zz__zz_stateReg_98_6 ? _zz__zz_stateReg_98_7 : _zz_stateReg_296)) ^ (_zz_stateReg_82[7] ? (_zz_stateReg_297 ^ _zz__zz_stateReg_98_8) : _zz_stateReg_297))) ^ (((_zz_stateReg_301[7] ? (_zz_stateReg_302 ^ _zz__zz_stateReg_98_9) : _zz_stateReg_302) ^ (_zz_stateReg_83[7] ? (_zz_stateReg_303 ^ _zz__zz_stateReg_98_10) : _zz_stateReg_303)) ^ _zz_stateReg_83));
    end
  end

  always @(*) begin
    _zz_stateReg_99 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_99 = _zz_stateReg_83;
    end else begin
      _zz_stateReg_99 = (((((_zz__zz_stateReg_99 ^ _zz__zz_stateReg_99_1) ^ _zz_stateReg_80) ^ ((_zz__zz_stateReg_99_2 ^ _zz__zz_stateReg_99_3) ^ _zz_stateReg_81)) ^ ((_zz_stateReg_321[7] ? (_zz_stateReg_322 ^ _zz__zz_stateReg_99_4) : _zz_stateReg_322) ^ _zz_stateReg_82)) ^ (((_zz_stateReg_326[7] ? (_zz_stateReg_327 ^ _zz__zz_stateReg_99_5) : _zz_stateReg_327) ^ (_zz_stateReg_329[7] ? (_zz_stateReg_330 ^ _zz__zz_stateReg_99_6) : _zz_stateReg_330)) ^ (_zz_stateReg_83[7] ? (_zz_stateReg_331 ^ 8'h1b) : _zz_stateReg_331)));
    end
  end

  always @(*) begin
    _zz_stateReg_100 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_100 = _zz_stateReg_84;
    end else begin
      _zz_stateReg_100 = (((((_zz__zz_stateReg_100 ^ _zz__zz_stateReg_100_1) ^ (_zz__zz_stateReg_100_2 ? _zz__zz_stateReg_100_3 : _zz_stateReg_340)) ^ ((_zz__zz_stateReg_100_4 ^ _zz__zz_stateReg_100_5) ^ _zz_stateReg_85)) ^ (((_zz__zz_stateReg_100_6 ? _zz__zz_stateReg_100_7 : _zz_stateReg_351) ^ (_zz__zz_stateReg_100_8 ? _zz__zz_stateReg_100_9 : _zz_stateReg_354)) ^ _zz_stateReg_86)) ^ ((_zz_stateReg_358[7] ? (_zz_stateReg_359 ^ 8'h1b) : _zz_stateReg_359) ^ _zz_stateReg_87));
    end
  end

  always @(*) begin
    _zz_stateReg_101 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_101 = _zz_stateReg_85;
    end else begin
      _zz_stateReg_101 = (((((_zz__zz_stateReg_101 ? _zz__zz_stateReg_101_1 : _zz_stateReg_364) ^ _zz_stateReg_84) ^ ((_zz__zz_stateReg_101_2 ^ _zz__zz_stateReg_101_3) ^ (_zz__zz_stateReg_101_4 ? _zz__zz_stateReg_101_5 : _zz_stateReg_373))) ^ (((_zz__zz_stateReg_101_6 ? _zz__zz_stateReg_101_7 : _zz_stateReg_378) ^ (_zz__zz_stateReg_101_8 ? _zz__zz_stateReg_101_9 : _zz_stateReg_379)) ^ _zz_stateReg_86)) ^ (((_zz_stateReg_383[7] ? (_zz_stateReg_384 ^ _zz__zz_stateReg_101_10) : _zz_stateReg_384) ^ (_zz_stateReg_386[7] ? (_zz_stateReg_387 ^ _zz__zz_stateReg_101_11) : _zz_stateReg_387)) ^ _zz_stateReg_87));
    end
  end

  always @(*) begin
    _zz_stateReg_102 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_102 = _zz_stateReg_86;
    end else begin
      _zz_stateReg_102 = (((((_zz__zz_stateReg_102 ^ _zz__zz_stateReg_102_1) ^ _zz_stateReg_84) ^ ((_zz__zz_stateReg_102_2 ? _zz__zz_stateReg_102_3 : _zz_stateReg_400) ^ _zz_stateReg_85)) ^ (((_zz__zz_stateReg_102_4 ? _zz__zz_stateReg_102_5 : _zz_stateReg_405) ^ (_zz__zz_stateReg_102_6 ? _zz__zz_stateReg_102_7 : _zz_stateReg_408)) ^ (_zz_stateReg_86[7] ? (_zz_stateReg_409 ^ _zz__zz_stateReg_102_8) : _zz_stateReg_409))) ^ (((_zz_stateReg_413[7] ? (_zz_stateReg_414 ^ _zz__zz_stateReg_102_9) : _zz_stateReg_414) ^ (_zz_stateReg_87[7] ? (_zz_stateReg_415 ^ _zz__zz_stateReg_102_10) : _zz_stateReg_415)) ^ _zz_stateReg_87));
    end
  end

  always @(*) begin
    _zz_stateReg_103 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_103 = _zz_stateReg_87;
    end else begin
      _zz_stateReg_103 = (((((_zz__zz_stateReg_103 ^ _zz__zz_stateReg_103_1) ^ _zz_stateReg_84) ^ ((_zz__zz_stateReg_103_2 ^ _zz__zz_stateReg_103_3) ^ _zz_stateReg_85)) ^ ((_zz_stateReg_433[7] ? (_zz_stateReg_434 ^ _zz__zz_stateReg_103_4) : _zz_stateReg_434) ^ _zz_stateReg_86)) ^ (((_zz_stateReg_438[7] ? (_zz_stateReg_439 ^ _zz__zz_stateReg_103_5) : _zz_stateReg_439) ^ (_zz_stateReg_441[7] ? (_zz_stateReg_442 ^ _zz__zz_stateReg_103_6) : _zz_stateReg_442)) ^ (_zz_stateReg_87[7] ? (_zz_stateReg_443 ^ 8'h1b) : _zz_stateReg_443)));
    end
  end

  always @(*) begin
    _zz_stateReg_104 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_104 = _zz_stateReg_88;
    end else begin
      _zz_stateReg_104 = (((((_zz__zz_stateReg_104 ^ _zz__zz_stateReg_104_1) ^ (_zz__zz_stateReg_104_2 ? _zz__zz_stateReg_104_3 : _zz_stateReg_452)) ^ ((_zz__zz_stateReg_104_4 ^ _zz__zz_stateReg_104_5) ^ _zz_stateReg_89)) ^ (((_zz__zz_stateReg_104_6 ? _zz__zz_stateReg_104_7 : _zz_stateReg_463) ^ (_zz__zz_stateReg_104_8 ? _zz__zz_stateReg_104_9 : _zz_stateReg_466)) ^ _zz_stateReg_90)) ^ ((_zz_stateReg_470[7] ? (_zz_stateReg_471 ^ 8'h1b) : _zz_stateReg_471) ^ _zz_stateReg_91));
    end
  end

  always @(*) begin
    _zz_stateReg_105 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_105 = _zz_stateReg_89;
    end else begin
      _zz_stateReg_105 = (((((_zz__zz_stateReg_105 ? _zz__zz_stateReg_105_1 : _zz_stateReg_476) ^ _zz_stateReg_88) ^ ((_zz__zz_stateReg_105_2 ^ _zz__zz_stateReg_105_3) ^ (_zz__zz_stateReg_105_4 ? _zz__zz_stateReg_105_5 : _zz_stateReg_485))) ^ (((_zz__zz_stateReg_105_6 ? _zz__zz_stateReg_105_7 : _zz_stateReg_490) ^ (_zz__zz_stateReg_105_8 ? _zz__zz_stateReg_105_9 : _zz_stateReg_491)) ^ _zz_stateReg_90)) ^ (((_zz_stateReg_495[7] ? (_zz_stateReg_496 ^ _zz__zz_stateReg_105_10) : _zz_stateReg_496) ^ (_zz_stateReg_498[7] ? (_zz_stateReg_499 ^ _zz__zz_stateReg_105_11) : _zz_stateReg_499)) ^ _zz_stateReg_91));
    end
  end

  always @(*) begin
    _zz_stateReg_106 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_106 = _zz_stateReg_90;
    end else begin
      _zz_stateReg_106 = (((((_zz__zz_stateReg_106 ^ _zz__zz_stateReg_106_1) ^ _zz_stateReg_88) ^ ((_zz__zz_stateReg_106_2 ? _zz__zz_stateReg_106_3 : _zz_stateReg_512) ^ _zz_stateReg_89)) ^ (((_zz__zz_stateReg_106_4 ? _zz__zz_stateReg_106_5 : _zz_stateReg_517) ^ (_zz__zz_stateReg_106_6 ? _zz__zz_stateReg_106_7 : _zz_stateReg_520)) ^ (_zz_stateReg_90[7] ? (_zz_stateReg_521 ^ _zz__zz_stateReg_106_8) : _zz_stateReg_521))) ^ (((_zz_stateReg_525[7] ? (_zz_stateReg_526 ^ _zz__zz_stateReg_106_9) : _zz_stateReg_526) ^ (_zz_stateReg_91[7] ? (_zz_stateReg_527 ^ _zz__zz_stateReg_106_10) : _zz_stateReg_527)) ^ _zz_stateReg_91));
    end
  end

  always @(*) begin
    _zz_stateReg_107 = 8'h0;
    if(when_AES128_l356) begin
      _zz_stateReg_107 = _zz_stateReg_91;
    end else begin
      _zz_stateReg_107 = (((((_zz__zz_stateReg_107 ^ _zz__zz_stateReg_107_1) ^ _zz_stateReg_88) ^ ((_zz__zz_stateReg_107_2 ^ _zz__zz_stateReg_107_3) ^ _zz_stateReg_89)) ^ ((_zz_stateReg_545[7] ? (_zz_stateReg_546 ^ _zz__zz_stateReg_107_4) : _zz_stateReg_546) ^ _zz_stateReg_90)) ^ (((_zz_stateReg_550[7] ? (_zz_stateReg_551 ^ _zz__zz_stateReg_107_5) : _zz_stateReg_551) ^ (_zz_stateReg_553[7] ? (_zz_stateReg_554 ^ _zz__zz_stateReg_107_6) : _zz_stateReg_554)) ^ (_zz_stateReg_91[7] ? (_zz_stateReg_555 ^ 8'h1b) : _zz_stateReg_555)));
    end
  end

  assign when_AES128_l356 = (rconCounter == 4'b0000);
  assign _zz_stateReg_108 = _zz__zz_stateReg_108[7 : 0];
  assign _zz_stateReg_109 = (_zz_stateReg_76[7] ? (_zz_stateReg_108 ^ 8'h1b) : _zz_stateReg_108);
  assign _zz_stateReg_110 = _zz__zz_stateReg_110[7 : 0];
  assign _zz_stateReg_111 = (_zz_stateReg_109[7] ? (_zz_stateReg_110 ^ 8'h1b) : _zz_stateReg_110);
  assign _zz_stateReg_112 = _zz__zz_stateReg_112[7 : 0];
  assign _zz_stateReg_113 = _zz__zz_stateReg_113[7 : 0];
  assign _zz_stateReg_114 = (_zz_stateReg_76[7] ? (_zz_stateReg_113 ^ 8'h1b) : _zz_stateReg_113);
  assign _zz_stateReg_115 = _zz__zz_stateReg_115[7 : 0];
  assign _zz_stateReg_116 = _zz__zz_stateReg_116[7 : 0];
  assign _zz_stateReg_117 = _zz__zz_stateReg_117[7 : 0];
  assign _zz_stateReg_118 = (_zz_stateReg_77[7] ? (_zz_stateReg_117 ^ 8'h1b) : _zz_stateReg_117);
  assign _zz_stateReg_119 = _zz__zz_stateReg_119[7 : 0];
  assign _zz_stateReg_120 = (_zz_stateReg_118[7] ? (_zz_stateReg_119 ^ 8'h1b) : _zz_stateReg_119);
  assign _zz_stateReg_121 = _zz__zz_stateReg_121[7 : 0];
  assign _zz_stateReg_122 = _zz__zz_stateReg_122[7 : 0];
  assign _zz_stateReg_123 = _zz__zz_stateReg_123[7 : 0];
  assign _zz_stateReg_124 = (_zz_stateReg_78[7] ? (_zz_stateReg_123 ^ 8'h1b) : _zz_stateReg_123);
  assign _zz_stateReg_125 = _zz__zz_stateReg_125[7 : 0];
  assign _zz_stateReg_126 = (_zz_stateReg_124[7] ? (_zz_stateReg_125 ^ 8'h1b) : _zz_stateReg_125);
  assign _zz_stateReg_127 = _zz__zz_stateReg_127[7 : 0];
  assign _zz_stateReg_128 = _zz__zz_stateReg_128[7 : 0];
  assign _zz_stateReg_129 = (_zz_stateReg_78[7] ? (_zz_stateReg_128 ^ 8'h1b) : _zz_stateReg_128);
  assign _zz_stateReg_130 = _zz__zz_stateReg_130[7 : 0];
  assign _zz_stateReg_131 = _zz__zz_stateReg_131[7 : 0];
  assign _zz_stateReg_132 = (_zz_stateReg_79[7] ? (_zz_stateReg_131 ^ 8'h1b) : _zz_stateReg_131);
  assign _zz_stateReg_133 = _zz__zz_stateReg_133[7 : 0];
  assign _zz_stateReg_134 = (_zz_stateReg_132[7] ? (_zz_stateReg_133 ^ 8'h1b) : _zz_stateReg_133);
  assign _zz_stateReg_135 = _zz__zz_stateReg_135[7 : 0];
  assign _zz_stateReg_136 = _zz__zz_stateReg_136[7 : 0];
  assign _zz_stateReg_137 = (_zz_stateReg_76[7] ? (_zz_stateReg_136 ^ 8'h1b) : _zz_stateReg_136);
  assign _zz_stateReg_138 = _zz__zz_stateReg_138[7 : 0];
  assign _zz_stateReg_139 = (_zz_stateReg_137[7] ? (_zz_stateReg_138 ^ 8'h1b) : _zz_stateReg_138);
  assign _zz_stateReg_140 = _zz__zz_stateReg_140[7 : 0];
  assign _zz_stateReg_141 = _zz__zz_stateReg_141[7 : 0];
  assign _zz_stateReg_142 = (_zz_stateReg_77[7] ? (_zz_stateReg_141 ^ 8'h1b) : _zz_stateReg_141);
  assign _zz_stateReg_143 = _zz__zz_stateReg_143[7 : 0];
  assign _zz_stateReg_144 = (_zz_stateReg_142[7] ? (_zz_stateReg_143 ^ 8'h1b) : _zz_stateReg_143);
  assign _zz_stateReg_145 = _zz__zz_stateReg_145[7 : 0];
  assign _zz_stateReg_146 = _zz__zz_stateReg_146[7 : 0];
  assign _zz_stateReg_147 = (_zz_stateReg_77[7] ? (_zz_stateReg_146 ^ 8'h1b) : _zz_stateReg_146);
  assign _zz_stateReg_148 = _zz__zz_stateReg_148[7 : 0];
  assign _zz_stateReg_149 = _zz__zz_stateReg_149[7 : 0];
  assign _zz_stateReg_150 = _zz__zz_stateReg_150[7 : 0];
  assign _zz_stateReg_151 = (_zz_stateReg_78[7] ? (_zz_stateReg_150 ^ 8'h1b) : _zz_stateReg_150);
  assign _zz_stateReg_152 = _zz__zz_stateReg_152[7 : 0];
  assign _zz_stateReg_153 = (_zz_stateReg_151[7] ? (_zz_stateReg_152 ^ 8'h1b) : _zz_stateReg_152);
  assign _zz_stateReg_154 = _zz__zz_stateReg_154[7 : 0];
  assign _zz_stateReg_155 = _zz__zz_stateReg_155[7 : 0];
  assign _zz_stateReg_156 = _zz__zz_stateReg_156[7 : 0];
  assign _zz_stateReg_157 = (_zz_stateReg_79[7] ? (_zz_stateReg_156 ^ 8'h1b) : _zz_stateReg_156);
  assign _zz_stateReg_158 = _zz__zz_stateReg_158[7 : 0];
  assign _zz_stateReg_159 = (_zz_stateReg_157[7] ? (_zz_stateReg_158 ^ 8'h1b) : _zz_stateReg_158);
  assign _zz_stateReg_160 = _zz__zz_stateReg_160[7 : 0];
  assign _zz_stateReg_161 = _zz__zz_stateReg_161[7 : 0];
  assign _zz_stateReg_162 = (_zz_stateReg_79[7] ? (_zz_stateReg_161 ^ 8'h1b) : _zz_stateReg_161);
  assign _zz_stateReg_163 = _zz__zz_stateReg_163[7 : 0];
  assign _zz_stateReg_164 = _zz__zz_stateReg_164[7 : 0];
  assign _zz_stateReg_165 = (_zz_stateReg_76[7] ? (_zz_stateReg_164 ^ 8'h1b) : _zz_stateReg_164);
  assign _zz_stateReg_166 = _zz__zz_stateReg_166[7 : 0];
  assign _zz_stateReg_167 = (_zz_stateReg_165[7] ? (_zz_stateReg_166 ^ 8'h1b) : _zz_stateReg_166);
  assign _zz_stateReg_168 = _zz__zz_stateReg_168[7 : 0];
  assign _zz_stateReg_169 = _zz__zz_stateReg_169[7 : 0];
  assign _zz_stateReg_170 = (_zz_stateReg_76[7] ? (_zz_stateReg_169 ^ 8'h1b) : _zz_stateReg_169);
  assign _zz_stateReg_171 = _zz__zz_stateReg_171[7 : 0];
  assign _zz_stateReg_172 = _zz__zz_stateReg_172[7 : 0];
  assign _zz_stateReg_173 = (_zz_stateReg_77[7] ? (_zz_stateReg_172 ^ 8'h1b) : _zz_stateReg_172);
  assign _zz_stateReg_174 = _zz__zz_stateReg_174[7 : 0];
  assign _zz_stateReg_175 = (_zz_stateReg_173[7] ? (_zz_stateReg_174 ^ 8'h1b) : _zz_stateReg_174);
  assign _zz_stateReg_176 = _zz__zz_stateReg_176[7 : 0];
  assign _zz_stateReg_177 = _zz__zz_stateReg_177[7 : 0];
  assign _zz_stateReg_178 = (_zz_stateReg_78[7] ? (_zz_stateReg_177 ^ 8'h1b) : _zz_stateReg_177);
  assign _zz_stateReg_179 = _zz__zz_stateReg_179[7 : 0];
  assign _zz_stateReg_180 = (_zz_stateReg_178[7] ? (_zz_stateReg_179 ^ 8'h1b) : _zz_stateReg_179);
  assign _zz_stateReg_181 = _zz__zz_stateReg_181[7 : 0];
  assign _zz_stateReg_182 = _zz__zz_stateReg_182[7 : 0];
  assign _zz_stateReg_183 = (_zz_stateReg_78[7] ? (_zz_stateReg_182 ^ 8'h1b) : _zz_stateReg_182);
  assign _zz_stateReg_184 = _zz__zz_stateReg_184[7 : 0];
  assign _zz_stateReg_185 = _zz__zz_stateReg_185[7 : 0];
  assign _zz_stateReg_186 = _zz__zz_stateReg_186[7 : 0];
  assign _zz_stateReg_187 = (_zz_stateReg_79[7] ? (_zz_stateReg_186 ^ 8'h1b) : _zz_stateReg_186);
  assign _zz_stateReg_188 = _zz__zz_stateReg_188[7 : 0];
  assign _zz_stateReg_189 = (_zz_stateReg_187[7] ? (_zz_stateReg_188 ^ 8'h1b) : _zz_stateReg_188);
  assign _zz_stateReg_190 = _zz__zz_stateReg_190[7 : 0];
  assign _zz_stateReg_191 = _zz__zz_stateReg_191[7 : 0];
  assign _zz_stateReg_192 = _zz__zz_stateReg_192[7 : 0];
  assign _zz_stateReg_193 = (_zz_stateReg_76[7] ? (_zz_stateReg_192 ^ 8'h1b) : _zz_stateReg_192);
  assign _zz_stateReg_194 = _zz__zz_stateReg_194[7 : 0];
  assign _zz_stateReg_195 = (_zz_stateReg_193[7] ? (_zz_stateReg_194 ^ 8'h1b) : _zz_stateReg_194);
  assign _zz_stateReg_196 = _zz__zz_stateReg_196[7 : 0];
  assign _zz_stateReg_197 = _zz__zz_stateReg_197[7 : 0];
  assign _zz_stateReg_198 = _zz__zz_stateReg_198[7 : 0];
  assign _zz_stateReg_199 = (_zz_stateReg_77[7] ? (_zz_stateReg_198 ^ 8'h1b) : _zz_stateReg_198);
  assign _zz_stateReg_200 = _zz__zz_stateReg_200[7 : 0];
  assign _zz_stateReg_201 = (_zz_stateReg_199[7] ? (_zz_stateReg_200 ^ 8'h1b) : _zz_stateReg_200);
  assign _zz_stateReg_202 = _zz__zz_stateReg_202[7 : 0];
  assign _zz_stateReg_203 = _zz__zz_stateReg_203[7 : 0];
  assign _zz_stateReg_204 = (_zz_stateReg_77[7] ? (_zz_stateReg_203 ^ 8'h1b) : _zz_stateReg_203);
  assign _zz_stateReg_205 = _zz__zz_stateReg_205[7 : 0];
  assign _zz_stateReg_206 = _zz__zz_stateReg_206[7 : 0];
  assign _zz_stateReg_207 = (_zz_stateReg_78[7] ? (_zz_stateReg_206 ^ 8'h1b) : _zz_stateReg_206);
  assign _zz_stateReg_208 = _zz__zz_stateReg_208[7 : 0];
  assign _zz_stateReg_209 = (_zz_stateReg_207[7] ? (_zz_stateReg_208 ^ 8'h1b) : _zz_stateReg_208);
  assign _zz_stateReg_210 = _zz__zz_stateReg_210[7 : 0];
  assign _zz_stateReg_211 = _zz__zz_stateReg_211[7 : 0];
  assign _zz_stateReg_212 = (_zz_stateReg_79[7] ? (_zz_stateReg_211 ^ 8'h1b) : _zz_stateReg_211);
  assign _zz_stateReg_213 = _zz__zz_stateReg_213[7 : 0];
  assign _zz_stateReg_214 = (_zz_stateReg_212[7] ? (_zz_stateReg_213 ^ 8'h1b) : _zz_stateReg_213);
  assign _zz_stateReg_215 = _zz__zz_stateReg_215[7 : 0];
  assign _zz_stateReg_216 = _zz__zz_stateReg_216[7 : 0];
  assign _zz_stateReg_217 = (_zz_stateReg_79[7] ? (_zz_stateReg_216 ^ 8'h1b) : _zz_stateReg_216);
  assign _zz_stateReg_218 = _zz__zz_stateReg_218[7 : 0];
  assign _zz_stateReg_219 = _zz__zz_stateReg_219[7 : 0];
  assign _zz_stateReg_220 = _zz__zz_stateReg_220[7 : 0];
  assign _zz_stateReg_221 = (_zz_stateReg_80[7] ? (_zz_stateReg_220 ^ 8'h1b) : _zz_stateReg_220);
  assign _zz_stateReg_222 = _zz__zz_stateReg_222[7 : 0];
  assign _zz_stateReg_223 = (_zz_stateReg_221[7] ? (_zz_stateReg_222 ^ 8'h1b) : _zz_stateReg_222);
  assign _zz_stateReg_224 = _zz__zz_stateReg_224[7 : 0];
  assign _zz_stateReg_225 = _zz__zz_stateReg_225[7 : 0];
  assign _zz_stateReg_226 = (_zz_stateReg_80[7] ? (_zz_stateReg_225 ^ 8'h1b) : _zz_stateReg_225);
  assign _zz_stateReg_227 = _zz__zz_stateReg_227[7 : 0];
  assign _zz_stateReg_228 = _zz__zz_stateReg_228[7 : 0];
  assign _zz_stateReg_229 = _zz__zz_stateReg_229[7 : 0];
  assign _zz_stateReg_230 = (_zz_stateReg_81[7] ? (_zz_stateReg_229 ^ 8'h1b) : _zz_stateReg_229);
  assign _zz_stateReg_231 = _zz__zz_stateReg_231[7 : 0];
  assign _zz_stateReg_232 = (_zz_stateReg_230[7] ? (_zz_stateReg_231 ^ 8'h1b) : _zz_stateReg_231);
  assign _zz_stateReg_233 = _zz__zz_stateReg_233[7 : 0];
  assign _zz_stateReg_234 = _zz__zz_stateReg_234[7 : 0];
  assign _zz_stateReg_235 = _zz__zz_stateReg_235[7 : 0];
  assign _zz_stateReg_236 = (_zz_stateReg_82[7] ? (_zz_stateReg_235 ^ 8'h1b) : _zz_stateReg_235);
  assign _zz_stateReg_237 = _zz__zz_stateReg_237[7 : 0];
  assign _zz_stateReg_238 = (_zz_stateReg_236[7] ? (_zz_stateReg_237 ^ 8'h1b) : _zz_stateReg_237);
  assign _zz_stateReg_239 = _zz__zz_stateReg_239[7 : 0];
  assign _zz_stateReg_240 = _zz__zz_stateReg_240[7 : 0];
  assign _zz_stateReg_241 = (_zz_stateReg_82[7] ? (_zz_stateReg_240 ^ 8'h1b) : _zz_stateReg_240);
  assign _zz_stateReg_242 = _zz__zz_stateReg_242[7 : 0];
  assign _zz_stateReg_243 = _zz__zz_stateReg_243[7 : 0];
  assign _zz_stateReg_244 = (_zz_stateReg_83[7] ? (_zz_stateReg_243 ^ 8'h1b) : _zz_stateReg_243);
  assign _zz_stateReg_245 = _zz__zz_stateReg_245[7 : 0];
  assign _zz_stateReg_246 = (_zz_stateReg_244[7] ? (_zz_stateReg_245 ^ 8'h1b) : _zz_stateReg_245);
  assign _zz_stateReg_247 = _zz__zz_stateReg_247[7 : 0];
  assign _zz_stateReg_248 = _zz__zz_stateReg_248[7 : 0];
  assign _zz_stateReg_249 = (_zz_stateReg_80[7] ? (_zz_stateReg_248 ^ 8'h1b) : _zz_stateReg_248);
  assign _zz_stateReg_250 = _zz__zz_stateReg_250[7 : 0];
  assign _zz_stateReg_251 = (_zz_stateReg_249[7] ? (_zz_stateReg_250 ^ 8'h1b) : _zz_stateReg_250);
  assign _zz_stateReg_252 = _zz__zz_stateReg_252[7 : 0];
  assign _zz_stateReg_253 = _zz__zz_stateReg_253[7 : 0];
  assign _zz_stateReg_254 = (_zz_stateReg_81[7] ? (_zz_stateReg_253 ^ 8'h1b) : _zz_stateReg_253);
  assign _zz_stateReg_255 = _zz__zz_stateReg_255[7 : 0];
  assign _zz_stateReg_256 = (_zz_stateReg_254[7] ? (_zz_stateReg_255 ^ 8'h1b) : _zz_stateReg_255);
  assign _zz_stateReg_257 = _zz__zz_stateReg_257[7 : 0];
  assign _zz_stateReg_258 = _zz__zz_stateReg_258[7 : 0];
  assign _zz_stateReg_259 = (_zz_stateReg_81[7] ? (_zz_stateReg_258 ^ 8'h1b) : _zz_stateReg_258);
  assign _zz_stateReg_260 = _zz__zz_stateReg_260[7 : 0];
  assign _zz_stateReg_261 = _zz__zz_stateReg_261[7 : 0];
  assign _zz_stateReg_262 = _zz__zz_stateReg_262[7 : 0];
  assign _zz_stateReg_263 = (_zz_stateReg_82[7] ? (_zz_stateReg_262 ^ 8'h1b) : _zz_stateReg_262);
  assign _zz_stateReg_264 = _zz__zz_stateReg_264[7 : 0];
  assign _zz_stateReg_265 = (_zz_stateReg_263[7] ? (_zz_stateReg_264 ^ 8'h1b) : _zz_stateReg_264);
  assign _zz_stateReg_266 = _zz__zz_stateReg_266[7 : 0];
  assign _zz_stateReg_267 = _zz__zz_stateReg_267[7 : 0];
  assign _zz_stateReg_268 = _zz__zz_stateReg_268[7 : 0];
  assign _zz_stateReg_269 = (_zz_stateReg_83[7] ? (_zz_stateReg_268 ^ 8'h1b) : _zz_stateReg_268);
  assign _zz_stateReg_270 = _zz__zz_stateReg_270[7 : 0];
  assign _zz_stateReg_271 = (_zz_stateReg_269[7] ? (_zz_stateReg_270 ^ 8'h1b) : _zz_stateReg_270);
  assign _zz_stateReg_272 = _zz__zz_stateReg_272[7 : 0];
  assign _zz_stateReg_273 = _zz__zz_stateReg_273[7 : 0];
  assign _zz_stateReg_274 = (_zz_stateReg_83[7] ? (_zz_stateReg_273 ^ 8'h1b) : _zz_stateReg_273);
  assign _zz_stateReg_275 = _zz__zz_stateReg_275[7 : 0];
  assign _zz_stateReg_276 = _zz__zz_stateReg_276[7 : 0];
  assign _zz_stateReg_277 = (_zz_stateReg_80[7] ? (_zz_stateReg_276 ^ 8'h1b) : _zz_stateReg_276);
  assign _zz_stateReg_278 = _zz__zz_stateReg_278[7 : 0];
  assign _zz_stateReg_279 = (_zz_stateReg_277[7] ? (_zz_stateReg_278 ^ 8'h1b) : _zz_stateReg_278);
  assign _zz_stateReg_280 = _zz__zz_stateReg_280[7 : 0];
  assign _zz_stateReg_281 = _zz__zz_stateReg_281[7 : 0];
  assign _zz_stateReg_282 = (_zz_stateReg_80[7] ? (_zz_stateReg_281 ^ 8'h1b) : _zz_stateReg_281);
  assign _zz_stateReg_283 = _zz__zz_stateReg_283[7 : 0];
  assign _zz_stateReg_284 = _zz__zz_stateReg_284[7 : 0];
  assign _zz_stateReg_285 = (_zz_stateReg_81[7] ? (_zz_stateReg_284 ^ 8'h1b) : _zz_stateReg_284);
  assign _zz_stateReg_286 = _zz__zz_stateReg_286[7 : 0];
  assign _zz_stateReg_287 = (_zz_stateReg_285[7] ? (_zz_stateReg_286 ^ 8'h1b) : _zz_stateReg_286);
  assign _zz_stateReg_288 = _zz__zz_stateReg_288[7 : 0];
  assign _zz_stateReg_289 = _zz__zz_stateReg_289[7 : 0];
  assign _zz_stateReg_290 = (_zz_stateReg_82[7] ? (_zz_stateReg_289 ^ 8'h1b) : _zz_stateReg_289);
  assign _zz_stateReg_291 = _zz__zz_stateReg_291[7 : 0];
  assign _zz_stateReg_292 = (_zz_stateReg_290[7] ? (_zz_stateReg_291 ^ 8'h1b) : _zz_stateReg_291);
  assign _zz_stateReg_293 = _zz__zz_stateReg_293[7 : 0];
  assign _zz_stateReg_294 = _zz__zz_stateReg_294[7 : 0];
  assign _zz_stateReg_295 = (_zz_stateReg_82[7] ? (_zz_stateReg_294 ^ 8'h1b) : _zz_stateReg_294);
  assign _zz_stateReg_296 = _zz__zz_stateReg_296[7 : 0];
  assign _zz_stateReg_297 = _zz__zz_stateReg_297[7 : 0];
  assign _zz_stateReg_298 = _zz__zz_stateReg_298[7 : 0];
  assign _zz_stateReg_299 = (_zz_stateReg_83[7] ? (_zz_stateReg_298 ^ 8'h1b) : _zz_stateReg_298);
  assign _zz_stateReg_300 = _zz__zz_stateReg_300[7 : 0];
  assign _zz_stateReg_301 = (_zz_stateReg_299[7] ? (_zz_stateReg_300 ^ 8'h1b) : _zz_stateReg_300);
  assign _zz_stateReg_302 = _zz__zz_stateReg_302[7 : 0];
  assign _zz_stateReg_303 = _zz__zz_stateReg_303[7 : 0];
  assign _zz_stateReg_304 = _zz__zz_stateReg_304[7 : 0];
  assign _zz_stateReg_305 = (_zz_stateReg_80[7] ? (_zz_stateReg_304 ^ 8'h1b) : _zz_stateReg_304);
  assign _zz_stateReg_306 = _zz__zz_stateReg_306[7 : 0];
  assign _zz_stateReg_307 = (_zz_stateReg_305[7] ? (_zz_stateReg_306 ^ 8'h1b) : _zz_stateReg_306);
  assign _zz_stateReg_308 = _zz__zz_stateReg_308[7 : 0];
  assign _zz_stateReg_309 = _zz__zz_stateReg_309[7 : 0];
  assign _zz_stateReg_310 = _zz__zz_stateReg_310[7 : 0];
  assign _zz_stateReg_311 = (_zz_stateReg_81[7] ? (_zz_stateReg_310 ^ 8'h1b) : _zz_stateReg_310);
  assign _zz_stateReg_312 = _zz__zz_stateReg_312[7 : 0];
  assign _zz_stateReg_313 = (_zz_stateReg_311[7] ? (_zz_stateReg_312 ^ 8'h1b) : _zz_stateReg_312);
  assign _zz_stateReg_314 = _zz__zz_stateReg_314[7 : 0];
  assign _zz_stateReg_315 = _zz__zz_stateReg_315[7 : 0];
  assign _zz_stateReg_316 = (_zz_stateReg_81[7] ? (_zz_stateReg_315 ^ 8'h1b) : _zz_stateReg_315);
  assign _zz_stateReg_317 = _zz__zz_stateReg_317[7 : 0];
  assign _zz_stateReg_318 = _zz__zz_stateReg_318[7 : 0];
  assign _zz_stateReg_319 = (_zz_stateReg_82[7] ? (_zz_stateReg_318 ^ 8'h1b) : _zz_stateReg_318);
  assign _zz_stateReg_320 = _zz__zz_stateReg_320[7 : 0];
  assign _zz_stateReg_321 = (_zz_stateReg_319[7] ? (_zz_stateReg_320 ^ 8'h1b) : _zz_stateReg_320);
  assign _zz_stateReg_322 = _zz__zz_stateReg_322[7 : 0];
  assign _zz_stateReg_323 = _zz__zz_stateReg_323[7 : 0];
  assign _zz_stateReg_324 = (_zz_stateReg_83[7] ? (_zz_stateReg_323 ^ 8'h1b) : _zz_stateReg_323);
  assign _zz_stateReg_325 = _zz__zz_stateReg_325[7 : 0];
  assign _zz_stateReg_326 = (_zz_stateReg_324[7] ? (_zz_stateReg_325 ^ 8'h1b) : _zz_stateReg_325);
  assign _zz_stateReg_327 = _zz__zz_stateReg_327[7 : 0];
  assign _zz_stateReg_328 = _zz__zz_stateReg_328[7 : 0];
  assign _zz_stateReg_329 = (_zz_stateReg_83[7] ? (_zz_stateReg_328 ^ 8'h1b) : _zz_stateReg_328);
  assign _zz_stateReg_330 = _zz__zz_stateReg_330[7 : 0];
  assign _zz_stateReg_331 = _zz__zz_stateReg_331[7 : 0];
  assign _zz_stateReg_332 = _zz__zz_stateReg_332[7 : 0];
  assign _zz_stateReg_333 = (_zz_stateReg_84[7] ? (_zz_stateReg_332 ^ 8'h1b) : _zz_stateReg_332);
  assign _zz_stateReg_334 = _zz__zz_stateReg_334[7 : 0];
  assign _zz_stateReg_335 = (_zz_stateReg_333[7] ? (_zz_stateReg_334 ^ 8'h1b) : _zz_stateReg_334);
  assign _zz_stateReg_336 = _zz__zz_stateReg_336[7 : 0];
  assign _zz_stateReg_337 = _zz__zz_stateReg_337[7 : 0];
  assign _zz_stateReg_338 = (_zz_stateReg_84[7] ? (_zz_stateReg_337 ^ 8'h1b) : _zz_stateReg_337);
  assign _zz_stateReg_339 = _zz__zz_stateReg_339[7 : 0];
  assign _zz_stateReg_340 = _zz__zz_stateReg_340[7 : 0];
  assign _zz_stateReg_341 = _zz__zz_stateReg_341[7 : 0];
  assign _zz_stateReg_342 = (_zz_stateReg_85[7] ? (_zz_stateReg_341 ^ 8'h1b) : _zz_stateReg_341);
  assign _zz_stateReg_343 = _zz__zz_stateReg_343[7 : 0];
  assign _zz_stateReg_344 = (_zz_stateReg_342[7] ? (_zz_stateReg_343 ^ 8'h1b) : _zz_stateReg_343);
  assign _zz_stateReg_345 = _zz__zz_stateReg_345[7 : 0];
  assign _zz_stateReg_346 = _zz__zz_stateReg_346[7 : 0];
  assign _zz_stateReg_347 = _zz__zz_stateReg_347[7 : 0];
  assign _zz_stateReg_348 = (_zz_stateReg_86[7] ? (_zz_stateReg_347 ^ 8'h1b) : _zz_stateReg_347);
  assign _zz_stateReg_349 = _zz__zz_stateReg_349[7 : 0];
  assign _zz_stateReg_350 = (_zz_stateReg_348[7] ? (_zz_stateReg_349 ^ 8'h1b) : _zz_stateReg_349);
  assign _zz_stateReg_351 = _zz__zz_stateReg_351[7 : 0];
  assign _zz_stateReg_352 = _zz__zz_stateReg_352[7 : 0];
  assign _zz_stateReg_353 = (_zz_stateReg_86[7] ? (_zz_stateReg_352 ^ 8'h1b) : _zz_stateReg_352);
  assign _zz_stateReg_354 = _zz__zz_stateReg_354[7 : 0];
  assign _zz_stateReg_355 = _zz__zz_stateReg_355[7 : 0];
  assign _zz_stateReg_356 = (_zz_stateReg_87[7] ? (_zz_stateReg_355 ^ 8'h1b) : _zz_stateReg_355);
  assign _zz_stateReg_357 = _zz__zz_stateReg_357[7 : 0];
  assign _zz_stateReg_358 = (_zz_stateReg_356[7] ? (_zz_stateReg_357 ^ 8'h1b) : _zz_stateReg_357);
  assign _zz_stateReg_359 = _zz__zz_stateReg_359[7 : 0];
  assign _zz_stateReg_360 = _zz__zz_stateReg_360[7 : 0];
  assign _zz_stateReg_361 = (_zz_stateReg_84[7] ? (_zz_stateReg_360 ^ 8'h1b) : _zz_stateReg_360);
  assign _zz_stateReg_362 = _zz__zz_stateReg_362[7 : 0];
  assign _zz_stateReg_363 = (_zz_stateReg_361[7] ? (_zz_stateReg_362 ^ 8'h1b) : _zz_stateReg_362);
  assign _zz_stateReg_364 = _zz__zz_stateReg_364[7 : 0];
  assign _zz_stateReg_365 = _zz__zz_stateReg_365[7 : 0];
  assign _zz_stateReg_366 = (_zz_stateReg_85[7] ? (_zz_stateReg_365 ^ 8'h1b) : _zz_stateReg_365);
  assign _zz_stateReg_367 = _zz__zz_stateReg_367[7 : 0];
  assign _zz_stateReg_368 = (_zz_stateReg_366[7] ? (_zz_stateReg_367 ^ 8'h1b) : _zz_stateReg_367);
  assign _zz_stateReg_369 = _zz__zz_stateReg_369[7 : 0];
  assign _zz_stateReg_370 = _zz__zz_stateReg_370[7 : 0];
  assign _zz_stateReg_371 = (_zz_stateReg_85[7] ? (_zz_stateReg_370 ^ 8'h1b) : _zz_stateReg_370);
  assign _zz_stateReg_372 = _zz__zz_stateReg_372[7 : 0];
  assign _zz_stateReg_373 = _zz__zz_stateReg_373[7 : 0];
  assign _zz_stateReg_374 = _zz__zz_stateReg_374[7 : 0];
  assign _zz_stateReg_375 = (_zz_stateReg_86[7] ? (_zz_stateReg_374 ^ 8'h1b) : _zz_stateReg_374);
  assign _zz_stateReg_376 = _zz__zz_stateReg_376[7 : 0];
  assign _zz_stateReg_377 = (_zz_stateReg_375[7] ? (_zz_stateReg_376 ^ 8'h1b) : _zz_stateReg_376);
  assign _zz_stateReg_378 = _zz__zz_stateReg_378[7 : 0];
  assign _zz_stateReg_379 = _zz__zz_stateReg_379[7 : 0];
  assign _zz_stateReg_380 = _zz__zz_stateReg_380[7 : 0];
  assign _zz_stateReg_381 = (_zz_stateReg_87[7] ? (_zz_stateReg_380 ^ 8'h1b) : _zz_stateReg_380);
  assign _zz_stateReg_382 = _zz__zz_stateReg_382[7 : 0];
  assign _zz_stateReg_383 = (_zz_stateReg_381[7] ? (_zz_stateReg_382 ^ 8'h1b) : _zz_stateReg_382);
  assign _zz_stateReg_384 = _zz__zz_stateReg_384[7 : 0];
  assign _zz_stateReg_385 = _zz__zz_stateReg_385[7 : 0];
  assign _zz_stateReg_386 = (_zz_stateReg_87[7] ? (_zz_stateReg_385 ^ 8'h1b) : _zz_stateReg_385);
  assign _zz_stateReg_387 = _zz__zz_stateReg_387[7 : 0];
  assign _zz_stateReg_388 = _zz__zz_stateReg_388[7 : 0];
  assign _zz_stateReg_389 = (_zz_stateReg_84[7] ? (_zz_stateReg_388 ^ 8'h1b) : _zz_stateReg_388);
  assign _zz_stateReg_390 = _zz__zz_stateReg_390[7 : 0];
  assign _zz_stateReg_391 = (_zz_stateReg_389[7] ? (_zz_stateReg_390 ^ 8'h1b) : _zz_stateReg_390);
  assign _zz_stateReg_392 = _zz__zz_stateReg_392[7 : 0];
  assign _zz_stateReg_393 = _zz__zz_stateReg_393[7 : 0];
  assign _zz_stateReg_394 = (_zz_stateReg_84[7] ? (_zz_stateReg_393 ^ 8'h1b) : _zz_stateReg_393);
  assign _zz_stateReg_395 = _zz__zz_stateReg_395[7 : 0];
  assign _zz_stateReg_396 = _zz__zz_stateReg_396[7 : 0];
  assign _zz_stateReg_397 = (_zz_stateReg_85[7] ? (_zz_stateReg_396 ^ 8'h1b) : _zz_stateReg_396);
  assign _zz_stateReg_398 = _zz__zz_stateReg_398[7 : 0];
  assign _zz_stateReg_399 = (_zz_stateReg_397[7] ? (_zz_stateReg_398 ^ 8'h1b) : _zz_stateReg_398);
  assign _zz_stateReg_400 = _zz__zz_stateReg_400[7 : 0];
  assign _zz_stateReg_401 = _zz__zz_stateReg_401[7 : 0];
  assign _zz_stateReg_402 = (_zz_stateReg_86[7] ? (_zz_stateReg_401 ^ 8'h1b) : _zz_stateReg_401);
  assign _zz_stateReg_403 = _zz__zz_stateReg_403[7 : 0];
  assign _zz_stateReg_404 = (_zz_stateReg_402[7] ? (_zz_stateReg_403 ^ 8'h1b) : _zz_stateReg_403);
  assign _zz_stateReg_405 = _zz__zz_stateReg_405[7 : 0];
  assign _zz_stateReg_406 = _zz__zz_stateReg_406[7 : 0];
  assign _zz_stateReg_407 = (_zz_stateReg_86[7] ? (_zz_stateReg_406 ^ 8'h1b) : _zz_stateReg_406);
  assign _zz_stateReg_408 = _zz__zz_stateReg_408[7 : 0];
  assign _zz_stateReg_409 = _zz__zz_stateReg_409[7 : 0];
  assign _zz_stateReg_410 = _zz__zz_stateReg_410[7 : 0];
  assign _zz_stateReg_411 = (_zz_stateReg_87[7] ? (_zz_stateReg_410 ^ 8'h1b) : _zz_stateReg_410);
  assign _zz_stateReg_412 = _zz__zz_stateReg_412[7 : 0];
  assign _zz_stateReg_413 = (_zz_stateReg_411[7] ? (_zz_stateReg_412 ^ 8'h1b) : _zz_stateReg_412);
  assign _zz_stateReg_414 = _zz__zz_stateReg_414[7 : 0];
  assign _zz_stateReg_415 = _zz__zz_stateReg_415[7 : 0];
  assign _zz_stateReg_416 = _zz__zz_stateReg_416[7 : 0];
  assign _zz_stateReg_417 = (_zz_stateReg_84[7] ? (_zz_stateReg_416 ^ 8'h1b) : _zz_stateReg_416);
  assign _zz_stateReg_418 = _zz__zz_stateReg_418[7 : 0];
  assign _zz_stateReg_419 = (_zz_stateReg_417[7] ? (_zz_stateReg_418 ^ 8'h1b) : _zz_stateReg_418);
  assign _zz_stateReg_420 = _zz__zz_stateReg_420[7 : 0];
  assign _zz_stateReg_421 = _zz__zz_stateReg_421[7 : 0];
  assign _zz_stateReg_422 = _zz__zz_stateReg_422[7 : 0];
  assign _zz_stateReg_423 = (_zz_stateReg_85[7] ? (_zz_stateReg_422 ^ 8'h1b) : _zz_stateReg_422);
  assign _zz_stateReg_424 = _zz__zz_stateReg_424[7 : 0];
  assign _zz_stateReg_425 = (_zz_stateReg_423[7] ? (_zz_stateReg_424 ^ 8'h1b) : _zz_stateReg_424);
  assign _zz_stateReg_426 = _zz__zz_stateReg_426[7 : 0];
  assign _zz_stateReg_427 = _zz__zz_stateReg_427[7 : 0];
  assign _zz_stateReg_428 = (_zz_stateReg_85[7] ? (_zz_stateReg_427 ^ 8'h1b) : _zz_stateReg_427);
  assign _zz_stateReg_429 = _zz__zz_stateReg_429[7 : 0];
  assign _zz_stateReg_430 = _zz__zz_stateReg_430[7 : 0];
  assign _zz_stateReg_431 = (_zz_stateReg_86[7] ? (_zz_stateReg_430 ^ 8'h1b) : _zz_stateReg_430);
  assign _zz_stateReg_432 = _zz__zz_stateReg_432[7 : 0];
  assign _zz_stateReg_433 = (_zz_stateReg_431[7] ? (_zz_stateReg_432 ^ 8'h1b) : _zz_stateReg_432);
  assign _zz_stateReg_434 = _zz__zz_stateReg_434[7 : 0];
  assign _zz_stateReg_435 = _zz__zz_stateReg_435[7 : 0];
  assign _zz_stateReg_436 = (_zz_stateReg_87[7] ? (_zz_stateReg_435 ^ 8'h1b) : _zz_stateReg_435);
  assign _zz_stateReg_437 = _zz__zz_stateReg_437[7 : 0];
  assign _zz_stateReg_438 = (_zz_stateReg_436[7] ? (_zz_stateReg_437 ^ 8'h1b) : _zz_stateReg_437);
  assign _zz_stateReg_439 = _zz__zz_stateReg_439[7 : 0];
  assign _zz_stateReg_440 = _zz__zz_stateReg_440[7 : 0];
  assign _zz_stateReg_441 = (_zz_stateReg_87[7] ? (_zz_stateReg_440 ^ 8'h1b) : _zz_stateReg_440);
  assign _zz_stateReg_442 = _zz__zz_stateReg_442[7 : 0];
  assign _zz_stateReg_443 = _zz__zz_stateReg_443[7 : 0];
  assign _zz_stateReg_444 = _zz__zz_stateReg_444[7 : 0];
  assign _zz_stateReg_445 = (_zz_stateReg_88[7] ? (_zz_stateReg_444 ^ 8'h1b) : _zz_stateReg_444);
  assign _zz_stateReg_446 = _zz__zz_stateReg_446[7 : 0];
  assign _zz_stateReg_447 = (_zz_stateReg_445[7] ? (_zz_stateReg_446 ^ 8'h1b) : _zz_stateReg_446);
  assign _zz_stateReg_448 = _zz__zz_stateReg_448[7 : 0];
  assign _zz_stateReg_449 = _zz__zz_stateReg_449[7 : 0];
  assign _zz_stateReg_450 = (_zz_stateReg_88[7] ? (_zz_stateReg_449 ^ 8'h1b) : _zz_stateReg_449);
  assign _zz_stateReg_451 = _zz__zz_stateReg_451[7 : 0];
  assign _zz_stateReg_452 = _zz__zz_stateReg_452[7 : 0];
  assign _zz_stateReg_453 = _zz__zz_stateReg_453[7 : 0];
  assign _zz_stateReg_454 = (_zz_stateReg_89[7] ? (_zz_stateReg_453 ^ 8'h1b) : _zz_stateReg_453);
  assign _zz_stateReg_455 = _zz__zz_stateReg_455[7 : 0];
  assign _zz_stateReg_456 = (_zz_stateReg_454[7] ? (_zz_stateReg_455 ^ 8'h1b) : _zz_stateReg_455);
  assign _zz_stateReg_457 = _zz__zz_stateReg_457[7 : 0];
  assign _zz_stateReg_458 = _zz__zz_stateReg_458[7 : 0];
  assign _zz_stateReg_459 = _zz__zz_stateReg_459[7 : 0];
  assign _zz_stateReg_460 = (_zz_stateReg_90[7] ? (_zz_stateReg_459 ^ 8'h1b) : _zz_stateReg_459);
  assign _zz_stateReg_461 = _zz__zz_stateReg_461[7 : 0];
  assign _zz_stateReg_462 = (_zz_stateReg_460[7] ? (_zz_stateReg_461 ^ 8'h1b) : _zz_stateReg_461);
  assign _zz_stateReg_463 = _zz__zz_stateReg_463[7 : 0];
  assign _zz_stateReg_464 = _zz__zz_stateReg_464[7 : 0];
  assign _zz_stateReg_465 = (_zz_stateReg_90[7] ? (_zz_stateReg_464 ^ 8'h1b) : _zz_stateReg_464);
  assign _zz_stateReg_466 = _zz__zz_stateReg_466[7 : 0];
  assign _zz_stateReg_467 = _zz__zz_stateReg_467[7 : 0];
  assign _zz_stateReg_468 = (_zz_stateReg_91[7] ? (_zz_stateReg_467 ^ 8'h1b) : _zz_stateReg_467);
  assign _zz_stateReg_469 = _zz__zz_stateReg_469[7 : 0];
  assign _zz_stateReg_470 = (_zz_stateReg_468[7] ? (_zz_stateReg_469 ^ 8'h1b) : _zz_stateReg_469);
  assign _zz_stateReg_471 = _zz__zz_stateReg_471[7 : 0];
  assign _zz_stateReg_472 = _zz__zz_stateReg_472[7 : 0];
  assign _zz_stateReg_473 = (_zz_stateReg_88[7] ? (_zz_stateReg_472 ^ 8'h1b) : _zz_stateReg_472);
  assign _zz_stateReg_474 = _zz__zz_stateReg_474[7 : 0];
  assign _zz_stateReg_475 = (_zz_stateReg_473[7] ? (_zz_stateReg_474 ^ 8'h1b) : _zz_stateReg_474);
  assign _zz_stateReg_476 = _zz__zz_stateReg_476[7 : 0];
  assign _zz_stateReg_477 = _zz__zz_stateReg_477[7 : 0];
  assign _zz_stateReg_478 = (_zz_stateReg_89[7] ? (_zz_stateReg_477 ^ 8'h1b) : _zz_stateReg_477);
  assign _zz_stateReg_479 = _zz__zz_stateReg_479[7 : 0];
  assign _zz_stateReg_480 = (_zz_stateReg_478[7] ? (_zz_stateReg_479 ^ 8'h1b) : _zz_stateReg_479);
  assign _zz_stateReg_481 = _zz__zz_stateReg_481[7 : 0];
  assign _zz_stateReg_482 = _zz__zz_stateReg_482[7 : 0];
  assign _zz_stateReg_483 = (_zz_stateReg_89[7] ? (_zz_stateReg_482 ^ 8'h1b) : _zz_stateReg_482);
  assign _zz_stateReg_484 = _zz__zz_stateReg_484[7 : 0];
  assign _zz_stateReg_485 = _zz__zz_stateReg_485[7 : 0];
  assign _zz_stateReg_486 = _zz__zz_stateReg_486[7 : 0];
  assign _zz_stateReg_487 = (_zz_stateReg_90[7] ? (_zz_stateReg_486 ^ 8'h1b) : _zz_stateReg_486);
  assign _zz_stateReg_488 = _zz__zz_stateReg_488[7 : 0];
  assign _zz_stateReg_489 = (_zz_stateReg_487[7] ? (_zz_stateReg_488 ^ 8'h1b) : _zz_stateReg_488);
  assign _zz_stateReg_490 = _zz__zz_stateReg_490[7 : 0];
  assign _zz_stateReg_491 = _zz__zz_stateReg_491[7 : 0];
  assign _zz_stateReg_492 = _zz__zz_stateReg_492[7 : 0];
  assign _zz_stateReg_493 = (_zz_stateReg_91[7] ? (_zz_stateReg_492 ^ 8'h1b) : _zz_stateReg_492);
  assign _zz_stateReg_494 = _zz__zz_stateReg_494[7 : 0];
  assign _zz_stateReg_495 = (_zz_stateReg_493[7] ? (_zz_stateReg_494 ^ 8'h1b) : _zz_stateReg_494);
  assign _zz_stateReg_496 = _zz__zz_stateReg_496[7 : 0];
  assign _zz_stateReg_497 = _zz__zz_stateReg_497[7 : 0];
  assign _zz_stateReg_498 = (_zz_stateReg_91[7] ? (_zz_stateReg_497 ^ 8'h1b) : _zz_stateReg_497);
  assign _zz_stateReg_499 = _zz__zz_stateReg_499[7 : 0];
  assign _zz_stateReg_500 = _zz__zz_stateReg_500[7 : 0];
  assign _zz_stateReg_501 = (_zz_stateReg_88[7] ? (_zz_stateReg_500 ^ 8'h1b) : _zz_stateReg_500);
  assign _zz_stateReg_502 = _zz__zz_stateReg_502[7 : 0];
  assign _zz_stateReg_503 = (_zz_stateReg_501[7] ? (_zz_stateReg_502 ^ 8'h1b) : _zz_stateReg_502);
  assign _zz_stateReg_504 = _zz__zz_stateReg_504[7 : 0];
  assign _zz_stateReg_505 = _zz__zz_stateReg_505[7 : 0];
  assign _zz_stateReg_506 = (_zz_stateReg_88[7] ? (_zz_stateReg_505 ^ 8'h1b) : _zz_stateReg_505);
  assign _zz_stateReg_507 = _zz__zz_stateReg_507[7 : 0];
  assign _zz_stateReg_508 = _zz__zz_stateReg_508[7 : 0];
  assign _zz_stateReg_509 = (_zz_stateReg_89[7] ? (_zz_stateReg_508 ^ 8'h1b) : _zz_stateReg_508);
  assign _zz_stateReg_510 = _zz__zz_stateReg_510[7 : 0];
  assign _zz_stateReg_511 = (_zz_stateReg_509[7] ? (_zz_stateReg_510 ^ 8'h1b) : _zz_stateReg_510);
  assign _zz_stateReg_512 = _zz__zz_stateReg_512[7 : 0];
  assign _zz_stateReg_513 = _zz__zz_stateReg_513[7 : 0];
  assign _zz_stateReg_514 = (_zz_stateReg_90[7] ? (_zz_stateReg_513 ^ 8'h1b) : _zz_stateReg_513);
  assign _zz_stateReg_515 = _zz__zz_stateReg_515[7 : 0];
  assign _zz_stateReg_516 = (_zz_stateReg_514[7] ? (_zz_stateReg_515 ^ 8'h1b) : _zz_stateReg_515);
  assign _zz_stateReg_517 = _zz__zz_stateReg_517[7 : 0];
  assign _zz_stateReg_518 = _zz__zz_stateReg_518[7 : 0];
  assign _zz_stateReg_519 = (_zz_stateReg_90[7] ? (_zz_stateReg_518 ^ 8'h1b) : _zz_stateReg_518);
  assign _zz_stateReg_520 = _zz__zz_stateReg_520[7 : 0];
  assign _zz_stateReg_521 = _zz__zz_stateReg_521[7 : 0];
  assign _zz_stateReg_522 = _zz__zz_stateReg_522[7 : 0];
  assign _zz_stateReg_523 = (_zz_stateReg_91[7] ? (_zz_stateReg_522 ^ 8'h1b) : _zz_stateReg_522);
  assign _zz_stateReg_524 = _zz__zz_stateReg_524[7 : 0];
  assign _zz_stateReg_525 = (_zz_stateReg_523[7] ? (_zz_stateReg_524 ^ 8'h1b) : _zz_stateReg_524);
  assign _zz_stateReg_526 = _zz__zz_stateReg_526[7 : 0];
  assign _zz_stateReg_527 = _zz__zz_stateReg_527[7 : 0];
  assign _zz_stateReg_528 = _zz__zz_stateReg_528[7 : 0];
  assign _zz_stateReg_529 = (_zz_stateReg_88[7] ? (_zz_stateReg_528 ^ 8'h1b) : _zz_stateReg_528);
  assign _zz_stateReg_530 = _zz__zz_stateReg_530[7 : 0];
  assign _zz_stateReg_531 = (_zz_stateReg_529[7] ? (_zz_stateReg_530 ^ 8'h1b) : _zz_stateReg_530);
  assign _zz_stateReg_532 = _zz__zz_stateReg_532[7 : 0];
  assign _zz_stateReg_533 = _zz__zz_stateReg_533[7 : 0];
  assign _zz_stateReg_534 = _zz__zz_stateReg_534[7 : 0];
  assign _zz_stateReg_535 = (_zz_stateReg_89[7] ? (_zz_stateReg_534 ^ 8'h1b) : _zz_stateReg_534);
  assign _zz_stateReg_536 = _zz__zz_stateReg_536[7 : 0];
  assign _zz_stateReg_537 = (_zz_stateReg_535[7] ? (_zz_stateReg_536 ^ 8'h1b) : _zz_stateReg_536);
  assign _zz_stateReg_538 = _zz__zz_stateReg_538[7 : 0];
  assign _zz_stateReg_539 = _zz__zz_stateReg_539[7 : 0];
  assign _zz_stateReg_540 = (_zz_stateReg_89[7] ? (_zz_stateReg_539 ^ 8'h1b) : _zz_stateReg_539);
  assign _zz_stateReg_541 = _zz__zz_stateReg_541[7 : 0];
  assign _zz_stateReg_542 = _zz__zz_stateReg_542[7 : 0];
  assign _zz_stateReg_543 = (_zz_stateReg_90[7] ? (_zz_stateReg_542 ^ 8'h1b) : _zz_stateReg_542);
  assign _zz_stateReg_544 = _zz__zz_stateReg_544[7 : 0];
  assign _zz_stateReg_545 = (_zz_stateReg_543[7] ? (_zz_stateReg_544 ^ 8'h1b) : _zz_stateReg_544);
  assign _zz_stateReg_546 = _zz__zz_stateReg_546[7 : 0];
  assign _zz_stateReg_547 = _zz__zz_stateReg_547[7 : 0];
  assign _zz_stateReg_548 = (_zz_stateReg_91[7] ? (_zz_stateReg_547 ^ 8'h1b) : _zz_stateReg_547);
  assign _zz_stateReg_549 = _zz__zz_stateReg_549[7 : 0];
  assign _zz_stateReg_550 = (_zz_stateReg_548[7] ? (_zz_stateReg_549 ^ 8'h1b) : _zz_stateReg_549);
  assign _zz_stateReg_551 = _zz__zz_stateReg_551[7 : 0];
  assign _zz_stateReg_552 = _zz__zz_stateReg_552[7 : 0];
  assign _zz_stateReg_553 = (_zz_stateReg_91[7] ? (_zz_stateReg_552 ^ 8'h1b) : _zz_stateReg_552);
  assign _zz_stateReg_554 = _zz__zz_stateReg_554[7 : 0];
  assign _zz_stateReg_555 = _zz__zz_stateReg_555[7 : 0];
  assign when_AES128_l383 = (roundCount == 4'b1010);
  assign when_AES128_l389 = (4'b0000 < rconCounter);
  assign when_AES128_l229 = (running && (! io_decrypt));
  assign when_AES128_l299 = (((! running) && (! precomputeRunning)) && io_decrypt);
  assign when_AES128_l324 = (running && io_decrypt);
  always @(posedge io_clk or posedge io_reset) begin
    if(io_reset) begin
      stateReg <= 128'h0;
      roundCount <= 4'b0000;
      running <= 1'b0;
      rconCounter <= 4'b0000;
      roundKeyReg_0 <= 32'h0;
      roundKeyReg_1 <= 32'h0;
      roundKeyReg_2 <= 32'h0;
      roundKeyReg_3 <= 32'h0;
      precomputeRunning <= 1'b0;
      precomputeCounter <= 4'b0000;
    end else begin
      if(when_AES128_l215) begin
        running <= 1'b1;
        stateReg <= {{{{{{_zz_stateReg_556,_zz_stateReg_568},_zz_stateReg_569},(_zz_stateReg_570 ^ _zz_stateReg_571)},(_zz_stateReg_572 ^ _zz_stateReg_3[23 : 16])},(io_dataIn[15 : 8] ^ _zz_stateReg_3[15 : 8])},(io_dataIn[7 : 0] ^ _zz_stateReg_3[7 : 0])};
        roundKeyReg_0 <= _zz_stateReg;
        roundKeyReg_1 <= _zz_stateReg_1;
        roundKeyReg_2 <= _zz_stateReg_2;
        roundKeyReg_3 <= _zz_stateReg_3;
        roundCount <= 4'b0000;
        rconCounter <= 4'b0000;
      end else begin
        if(when_AES128_l229) begin
          stateReg <= (_zz_stateReg_68 ^ _zz_stateReg_69);
          roundKeyReg_0 <= _zz_roundKeyReg_0_2;
          roundKeyReg_1 <= _zz_roundKeyReg_1;
          roundKeyReg_2 <= _zz_roundKeyReg_2;
          roundKeyReg_3 <= _zz_roundKeyReg_3;
          if(when_AES128_l291) begin
            running <= 1'b0;
          end else begin
            roundCount <= (roundCount + 4'b0001);
            if(when_AES128_l297) begin
              rconCounter <= (rconCounter + 4'b0001);
            end
          end
        end else begin
          if(when_AES128_l299) begin
            roundKeyReg_0 <= io_key[127 : 96];
            roundKeyReg_1 <= io_key[95 : 64];
            roundKeyReg_2 <= io_key[63 : 32];
            roundKeyReg_3 <= io_key[31 : 0];
            precomputeRunning <= 1'b1;
            precomputeCounter <= 4'b0000;
            rconCounter <= 4'b0000;
          end else begin
            if(precomputeRunning) begin
              roundKeyReg_0 <= _zz_stateReg_71;
              roundKeyReg_1 <= _zz_stateReg_72;
              roundKeyReg_2 <= _zz_stateReg_73;
              roundKeyReg_3 <= _zz_stateReg_74;
              precomputeCounter <= (precomputeCounter + 4'b0001);
              if(when_AES128_l313) begin
                precomputeRunning <= 1'b0;
                roundKeyReg_0 <= _zz_stateReg_71;
                roundKeyReg_1 <= _zz_stateReg_72;
                roundKeyReg_2 <= _zz_stateReg_73;
                roundKeyReg_3 <= _zz_stateReg_74;
                stateReg <= (io_dataIn ^ {{{{{{{{{_zz_stateReg_573,_zz_stateReg_574},_zz_stateReg_575},_zz_stateReg_73[23 : 16]},_zz_stateReg_73[15 : 8]},_zz_stateReg_73[7 : 0]},_zz_stateReg_74[31 : 24]},_zz_stateReg_74[23 : 16]},_zz_stateReg_74[15 : 8]},_zz_stateReg_74[7 : 0]});
                running <= 1'b1;
                roundCount <= 4'b0000;
                rconCounter <= 4'b1001;
              end
            end else begin
              if(when_AES128_l324) begin
                stateReg <= {{{{{{{{{{{_zz_stateReg_576,_zz_stateReg_577},_zz_stateReg_98},_zz_stateReg_99},_zz_stateReg_100},_zz_stateReg_101},_zz_stateReg_102},_zz_stateReg_103},_zz_stateReg_104},_zz_stateReg_105},_zz_stateReg_106},_zz_stateReg_107};
                roundKeyReg_0 <= _zz_roundKeyReg_0_4;
                roundKeyReg_1 <= _zz_roundKeyReg_1_1;
                roundKeyReg_2 <= _zz_roundKeyReg_2_1;
                roundKeyReg_3 <= _zz_roundKeyReg_3_1;
                if(when_AES128_l383) begin
                  running <= 1'b0;
                end else begin
                  roundCount <= (roundCount + 4'b0001);
                  if(when_AES128_l389) begin
                    rconCounter <= (rconCounter - 4'b0001);
                  end
                end
              end
            end
          end
        end
      end
    end
  end


endmodule
