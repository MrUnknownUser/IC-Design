// Generator : SpinalHDL v1.12.3    git head : 591e64062329e5e2e2b81f4d52422948053edb97
// Component : AesIterative
// Git hash  : c3e1a8c70c77e783c38c8c9886fb00a7b62a4b97

`timescale 1ns/1ps

module AesIterative (
  input  wire          io_start,
  input  wire [127:0]  io_key,
  input  wire [127:0]  io_dataIn,
  output reg  [127:0]  io_dataOut,
  output wire          io_busy,
  output reg           io_done,
  input  wire          clk,
  input  wire          reset
);

  wire       [79:0]   _zz_stateReg_70;
  wire       [39:0]   _zz_stateReg_71;
  wire       [7:0]    _zz_stateReg_72;
  wire       [7:0]    _zz_stateReg_73;
  wire       [7:0]    _zz_stateReg_74;
  wire       [7:0]    _zz_stateReg_75;
  wire       [7:0]    _zz_stateReg_76;
  wire       [7:0]    _zz_stateReg_77;
  wire       [7:0]    _zz_stateReg_78;
  wire       [7:0]    _zz_stateReg_79;
  wire       [7:0]    _zz_stateReg_80;
  wire       [7:0]    _zz_stateReg_81;
  wire       [7:0]    _zz_stateReg_82;
  wire       [7:0]    _zz_stateReg_83;
  wire       [7:0]    _zz_stateReg_84;
  wire       [7:0]    _zz_stateReg_85;
  wire       [7:0]    _zz_stateReg_86;
  reg        [7:0]    _zz__zz_stateReg_4;
  wire       [7:0]    _zz__zz_stateReg_4_1;
  reg        [7:0]    _zz__zz_stateReg_8;
  wire       [7:0]    _zz__zz_stateReg_8_1;
  reg        [7:0]    _zz__zz_stateReg_12;
  wire       [7:0]    _zz__zz_stateReg_12_1;
  reg        [7:0]    _zz__zz_stateReg_16;
  wire       [7:0]    _zz__zz_stateReg_16_1;
  reg        [7:0]    _zz__zz_stateReg_5;
  wire       [7:0]    _zz__zz_stateReg_5_1;
  reg        [7:0]    _zz__zz_stateReg_9;
  wire       [7:0]    _zz__zz_stateReg_9_1;
  reg        [7:0]    _zz__zz_stateReg_13;
  wire       [7:0]    _zz__zz_stateReg_13_1;
  reg        [7:0]    _zz__zz_stateReg_17;
  wire       [7:0]    _zz__zz_stateReg_17_1;
  reg        [7:0]    _zz__zz_stateReg_6;
  wire       [7:0]    _zz__zz_stateReg_6_1;
  reg        [7:0]    _zz__zz_stateReg_10;
  wire       [7:0]    _zz__zz_stateReg_10_1;
  reg        [7:0]    _zz__zz_stateReg_14;
  wire       [7:0]    _zz__zz_stateReg_14_1;
  reg        [7:0]    _zz__zz_stateReg_18;
  wire       [7:0]    _zz__zz_stateReg_18_1;
  reg        [7:0]    _zz__zz_stateReg_7;
  wire       [7:0]    _zz__zz_stateReg_7_1;
  reg        [7:0]    _zz__zz_stateReg_11;
  wire       [7:0]    _zz__zz_stateReg_11_1;
  reg        [7:0]    _zz__zz_stateReg_15;
  wire       [7:0]    _zz__zz_stateReg_15_1;
  reg        [7:0]    _zz__zz_stateReg_19;
  wire       [7:0]    _zz__zz_stateReg_19_1;
  wire       [8:0]    _zz__zz_stateReg_36;
  wire       [8:0]    _zz__zz_stateReg_37;
  wire       [8:0]    _zz__zz_stateReg_38;
  wire       [8:0]    _zz__zz_stateReg_39;
  wire       [8:0]    _zz__zz_stateReg_40;
  wire       [8:0]    _zz__zz_stateReg_41;
  wire       [8:0]    _zz__zz_stateReg_42;
  wire       [8:0]    _zz__zz_stateReg_43;
  wire       [8:0]    _zz__zz_stateReg_44;
  wire       [8:0]    _zz__zz_stateReg_45;
  wire       [8:0]    _zz__zz_stateReg_46;
  wire       [8:0]    _zz__zz_stateReg_47;
  wire       [8:0]    _zz__zz_stateReg_48;
  wire       [8:0]    _zz__zz_stateReg_49;
  wire       [8:0]    _zz__zz_stateReg_50;
  wire       [8:0]    _zz__zz_stateReg_51;
  wire       [8:0]    _zz__zz_stateReg_52;
  wire       [8:0]    _zz__zz_stateReg_53;
  wire       [8:0]    _zz__zz_stateReg_54;
  wire       [8:0]    _zz__zz_stateReg_55;
  wire       [8:0]    _zz__zz_stateReg_56;
  wire       [8:0]    _zz__zz_stateReg_57;
  wire       [8:0]    _zz__zz_stateReg_58;
  wire       [8:0]    _zz__zz_stateReg_59;
  wire       [8:0]    _zz__zz_stateReg_60;
  wire       [8:0]    _zz__zz_stateReg_61;
  wire       [8:0]    _zz__zz_stateReg_62;
  wire       [8:0]    _zz__zz_stateReg_63;
  wire       [8:0]    _zz__zz_stateReg_64;
  wire       [8:0]    _zz__zz_stateReg_65;
  wire       [8:0]    _zz__zz_stateReg_66;
  wire       [8:0]    _zz__zz_stateReg_67;
  wire       [39:0]   _zz__zz_stateReg_68;
  wire       [7:0]    _zz__zz_stateReg_68_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0_1;
  wire       [7:0]    _zz__zz_roundKeyReg_0_1_1;
  reg        [7:0]    _zz__zz_roundKeyReg_0_1_2;
  wire       [7:0]    _zz__zz_roundKeyReg_0_1_3;
  reg        [7:0]    _zz__zz_roundKeyReg_0_1_4;
  wire       [7:0]    _zz__zz_roundKeyReg_0_1_5;
  reg        [7:0]    _zz__zz_roundKeyReg_0_1_6;
  wire       [7:0]    _zz__zz_roundKeyReg_0_1_7;
  reg        [7:0]    _zz__zz_roundKeyReg_0_1_8;
  wire       [55:0]   _zz__zz_stateReg_69;
  wire       [7:0]    _zz__zz_stateReg_69_1;
  wire       [7:0]    _zz__zz_stateReg_69_2;
  wire       [7:0]    sboxRom_0;
  wire       [7:0]    sboxRom_1;
  wire       [7:0]    sboxRom_2;
  wire       [7:0]    sboxRom_3;
  wire       [7:0]    sboxRom_4;
  wire       [7:0]    sboxRom_5;
  wire       [7:0]    sboxRom_6;
  wire       [7:0]    sboxRom_7;
  wire       [7:0]    sboxRom_8;
  wire       [7:0]    sboxRom_9;
  wire       [7:0]    sboxRom_10;
  wire       [7:0]    sboxRom_11;
  wire       [7:0]    sboxRom_12;
  wire       [7:0]    sboxRom_13;
  wire       [7:0]    sboxRom_14;
  wire       [7:0]    sboxRom_15;
  wire       [7:0]    sboxRom_16;
  wire       [7:0]    sboxRom_17;
  wire       [7:0]    sboxRom_18;
  wire       [7:0]    sboxRom_19;
  wire       [7:0]    sboxRom_20;
  wire       [7:0]    sboxRom_21;
  wire       [7:0]    sboxRom_22;
  wire       [7:0]    sboxRom_23;
  wire       [7:0]    sboxRom_24;
  wire       [7:0]    sboxRom_25;
  wire       [7:0]    sboxRom_26;
  wire       [7:0]    sboxRom_27;
  wire       [7:0]    sboxRom_28;
  wire       [7:0]    sboxRom_29;
  wire       [7:0]    sboxRom_30;
  wire       [7:0]    sboxRom_31;
  wire       [7:0]    sboxRom_32;
  wire       [7:0]    sboxRom_33;
  wire       [7:0]    sboxRom_34;
  wire       [7:0]    sboxRom_35;
  wire       [7:0]    sboxRom_36;
  wire       [7:0]    sboxRom_37;
  wire       [7:0]    sboxRom_38;
  wire       [7:0]    sboxRom_39;
  wire       [7:0]    sboxRom_40;
  wire       [7:0]    sboxRom_41;
  wire       [7:0]    sboxRom_42;
  wire       [7:0]    sboxRom_43;
  wire       [7:0]    sboxRom_44;
  wire       [7:0]    sboxRom_45;
  wire       [7:0]    sboxRom_46;
  wire       [7:0]    sboxRom_47;
  wire       [7:0]    sboxRom_48;
  wire       [7:0]    sboxRom_49;
  wire       [7:0]    sboxRom_50;
  wire       [7:0]    sboxRom_51;
  wire       [7:0]    sboxRom_52;
  wire       [7:0]    sboxRom_53;
  wire       [7:0]    sboxRom_54;
  wire       [7:0]    sboxRom_55;
  wire       [7:0]    sboxRom_56;
  wire       [7:0]    sboxRom_57;
  wire       [7:0]    sboxRom_58;
  wire       [7:0]    sboxRom_59;
  wire       [7:0]    sboxRom_60;
  wire       [7:0]    sboxRom_61;
  wire       [7:0]    sboxRom_62;
  wire       [7:0]    sboxRom_63;
  wire       [7:0]    sboxRom_64;
  wire       [7:0]    sboxRom_65;
  wire       [7:0]    sboxRom_66;
  wire       [7:0]    sboxRom_67;
  wire       [7:0]    sboxRom_68;
  wire       [7:0]    sboxRom_69;
  wire       [7:0]    sboxRom_70;
  wire       [7:0]    sboxRom_71;
  wire       [7:0]    sboxRom_72;
  wire       [7:0]    sboxRom_73;
  wire       [7:0]    sboxRom_74;
  wire       [7:0]    sboxRom_75;
  wire       [7:0]    sboxRom_76;
  wire       [7:0]    sboxRom_77;
  wire       [7:0]    sboxRom_78;
  wire       [7:0]    sboxRom_79;
  wire       [7:0]    sboxRom_80;
  wire       [7:0]    sboxRom_81;
  wire       [7:0]    sboxRom_82;
  wire       [7:0]    sboxRom_83;
  wire       [7:0]    sboxRom_84;
  wire       [7:0]    sboxRom_85;
  wire       [7:0]    sboxRom_86;
  wire       [7:0]    sboxRom_87;
  wire       [7:0]    sboxRom_88;
  wire       [7:0]    sboxRom_89;
  wire       [7:0]    sboxRom_90;
  wire       [7:0]    sboxRom_91;
  wire       [7:0]    sboxRom_92;
  wire       [7:0]    sboxRom_93;
  wire       [7:0]    sboxRom_94;
  wire       [7:0]    sboxRom_95;
  wire       [7:0]    sboxRom_96;
  wire       [7:0]    sboxRom_97;
  wire       [7:0]    sboxRom_98;
  wire       [7:0]    sboxRom_99;
  wire       [7:0]    sboxRom_100;
  wire       [7:0]    sboxRom_101;
  wire       [7:0]    sboxRom_102;
  wire       [7:0]    sboxRom_103;
  wire       [7:0]    sboxRom_104;
  wire       [7:0]    sboxRom_105;
  wire       [7:0]    sboxRom_106;
  wire       [7:0]    sboxRom_107;
  wire       [7:0]    sboxRom_108;
  wire       [7:0]    sboxRom_109;
  wire       [7:0]    sboxRom_110;
  wire       [7:0]    sboxRom_111;
  wire       [7:0]    sboxRom_112;
  wire       [7:0]    sboxRom_113;
  wire       [7:0]    sboxRom_114;
  wire       [7:0]    sboxRom_115;
  wire       [7:0]    sboxRom_116;
  wire       [7:0]    sboxRom_117;
  wire       [7:0]    sboxRom_118;
  wire       [7:0]    sboxRom_119;
  wire       [7:0]    sboxRom_120;
  wire       [7:0]    sboxRom_121;
  wire       [7:0]    sboxRom_122;
  wire       [7:0]    sboxRom_123;
  wire       [7:0]    sboxRom_124;
  wire       [7:0]    sboxRom_125;
  wire       [7:0]    sboxRom_126;
  wire       [7:0]    sboxRom_127;
  wire       [7:0]    sboxRom_128;
  wire       [7:0]    sboxRom_129;
  wire       [7:0]    sboxRom_130;
  wire       [7:0]    sboxRom_131;
  wire       [7:0]    sboxRom_132;
  wire       [7:0]    sboxRom_133;
  wire       [7:0]    sboxRom_134;
  wire       [7:0]    sboxRom_135;
  wire       [7:0]    sboxRom_136;
  wire       [7:0]    sboxRom_137;
  wire       [7:0]    sboxRom_138;
  wire       [7:0]    sboxRom_139;
  wire       [7:0]    sboxRom_140;
  wire       [7:0]    sboxRom_141;
  wire       [7:0]    sboxRom_142;
  wire       [7:0]    sboxRom_143;
  wire       [7:0]    sboxRom_144;
  wire       [7:0]    sboxRom_145;
  wire       [7:0]    sboxRom_146;
  wire       [7:0]    sboxRom_147;
  wire       [7:0]    sboxRom_148;
  wire       [7:0]    sboxRom_149;
  wire       [7:0]    sboxRom_150;
  wire       [7:0]    sboxRom_151;
  wire       [7:0]    sboxRom_152;
  wire       [7:0]    sboxRom_153;
  wire       [7:0]    sboxRom_154;
  wire       [7:0]    sboxRom_155;
  wire       [7:0]    sboxRom_156;
  wire       [7:0]    sboxRom_157;
  wire       [7:0]    sboxRom_158;
  wire       [7:0]    sboxRom_159;
  wire       [7:0]    sboxRom_160;
  wire       [7:0]    sboxRom_161;
  wire       [7:0]    sboxRom_162;
  wire       [7:0]    sboxRom_163;
  wire       [7:0]    sboxRom_164;
  wire       [7:0]    sboxRom_165;
  wire       [7:0]    sboxRom_166;
  wire       [7:0]    sboxRom_167;
  wire       [7:0]    sboxRom_168;
  wire       [7:0]    sboxRom_169;
  wire       [7:0]    sboxRom_170;
  wire       [7:0]    sboxRom_171;
  wire       [7:0]    sboxRom_172;
  wire       [7:0]    sboxRom_173;
  wire       [7:0]    sboxRom_174;
  wire       [7:0]    sboxRom_175;
  wire       [7:0]    sboxRom_176;
  wire       [7:0]    sboxRom_177;
  wire       [7:0]    sboxRom_178;
  wire       [7:0]    sboxRom_179;
  wire       [7:0]    sboxRom_180;
  wire       [7:0]    sboxRom_181;
  wire       [7:0]    sboxRom_182;
  wire       [7:0]    sboxRom_183;
  wire       [7:0]    sboxRom_184;
  wire       [7:0]    sboxRom_185;
  wire       [7:0]    sboxRom_186;
  wire       [7:0]    sboxRom_187;
  wire       [7:0]    sboxRom_188;
  wire       [7:0]    sboxRom_189;
  wire       [7:0]    sboxRom_190;
  wire       [7:0]    sboxRom_191;
  wire       [7:0]    sboxRom_192;
  wire       [7:0]    sboxRom_193;
  wire       [7:0]    sboxRom_194;
  wire       [7:0]    sboxRom_195;
  wire       [7:0]    sboxRom_196;
  wire       [7:0]    sboxRom_197;
  wire       [7:0]    sboxRom_198;
  wire       [7:0]    sboxRom_199;
  wire       [7:0]    sboxRom_200;
  wire       [7:0]    sboxRom_201;
  wire       [7:0]    sboxRom_202;
  wire       [7:0]    sboxRom_203;
  wire       [7:0]    sboxRom_204;
  wire       [7:0]    sboxRom_205;
  wire       [7:0]    sboxRom_206;
  wire       [7:0]    sboxRom_207;
  wire       [7:0]    sboxRom_208;
  wire       [7:0]    sboxRom_209;
  wire       [7:0]    sboxRom_210;
  wire       [7:0]    sboxRom_211;
  wire       [7:0]    sboxRom_212;
  wire       [7:0]    sboxRom_213;
  wire       [7:0]    sboxRom_214;
  wire       [7:0]    sboxRom_215;
  wire       [7:0]    sboxRom_216;
  wire       [7:0]    sboxRom_217;
  wire       [7:0]    sboxRom_218;
  wire       [7:0]    sboxRom_219;
  wire       [7:0]    sboxRom_220;
  wire       [7:0]    sboxRom_221;
  wire       [7:0]    sboxRom_222;
  wire       [7:0]    sboxRom_223;
  wire       [7:0]    sboxRom_224;
  wire       [7:0]    sboxRom_225;
  wire       [7:0]    sboxRom_226;
  wire       [7:0]    sboxRom_227;
  wire       [7:0]    sboxRom_228;
  wire       [7:0]    sboxRom_229;
  wire       [7:0]    sboxRom_230;
  wire       [7:0]    sboxRom_231;
  wire       [7:0]    sboxRom_232;
  wire       [7:0]    sboxRom_233;
  wire       [7:0]    sboxRom_234;
  wire       [7:0]    sboxRom_235;
  wire       [7:0]    sboxRom_236;
  wire       [7:0]    sboxRom_237;
  wire       [7:0]    sboxRom_238;
  wire       [7:0]    sboxRom_239;
  wire       [7:0]    sboxRom_240;
  wire       [7:0]    sboxRom_241;
  wire       [7:0]    sboxRom_242;
  wire       [7:0]    sboxRom_243;
  wire       [7:0]    sboxRom_244;
  wire       [7:0]    sboxRom_245;
  wire       [7:0]    sboxRom_246;
  wire       [7:0]    sboxRom_247;
  wire       [7:0]    sboxRom_248;
  wire       [7:0]    sboxRom_249;
  wire       [7:0]    sboxRom_250;
  wire       [7:0]    sboxRom_251;
  wire       [7:0]    sboxRom_252;
  wire       [7:0]    sboxRom_253;
  wire       [7:0]    sboxRom_254;
  wire       [7:0]    sboxRom_255;
  wire       [7:0]    rcon_0;
  wire       [7:0]    rcon_1;
  wire       [7:0]    rcon_2;
  wire       [7:0]    rcon_3;
  wire       [7:0]    rcon_4;
  wire       [7:0]    rcon_5;
  wire       [7:0]    rcon_6;
  wire       [7:0]    rcon_7;
  wire       [7:0]    rcon_8;
  wire       [7:0]    rcon_9;
  reg        [127:0]  stateReg;
  reg        [31:0]   roundKeyReg_0;
  reg        [31:0]   roundKeyReg_1;
  reg        [31:0]   roundKeyReg_2;
  reg        [31:0]   roundKeyReg_3;
  reg        [3:0]    roundCount;
  reg                 running;
  reg        [3:0]    rconCounter;
  reg        [127:0]  newStateComb;
  reg        [127:0]  rkBitsUsedComb;
  wire                when_AES128_l150;
  wire       [31:0]   _zz_stateReg;
  wire       [31:0]   _zz_stateReg_1;
  wire       [31:0]   _zz_stateReg_2;
  wire       [31:0]   _zz_stateReg_3;
  wire       [7:0]    _zz_stateReg_4;
  wire       [7:0]    _zz_stateReg_5;
  wire       [7:0]    _zz_stateReg_6;
  wire       [7:0]    _zz_stateReg_7;
  wire       [7:0]    _zz_stateReg_8;
  wire       [7:0]    _zz_stateReg_9;
  wire       [7:0]    _zz_stateReg_10;
  wire       [7:0]    _zz_stateReg_11;
  wire       [7:0]    _zz_stateReg_12;
  wire       [7:0]    _zz_stateReg_13;
  wire       [7:0]    _zz_stateReg_14;
  wire       [7:0]    _zz_stateReg_15;
  wire       [7:0]    _zz_stateReg_16;
  wire       [7:0]    _zz_stateReg_17;
  wire       [7:0]    _zz_stateReg_18;
  wire       [7:0]    _zz_stateReg_19;
  reg        [7:0]    _zz_stateReg_20;
  reg        [7:0]    _zz_stateReg_21;
  reg        [7:0]    _zz_stateReg_22;
  reg        [7:0]    _zz_stateReg_23;
  reg        [7:0]    _zz_stateReg_24;
  reg        [7:0]    _zz_stateReg_25;
  reg        [7:0]    _zz_stateReg_26;
  reg        [7:0]    _zz_stateReg_27;
  reg        [7:0]    _zz_stateReg_28;
  reg        [7:0]    _zz_stateReg_29;
  reg        [7:0]    _zz_stateReg_30;
  reg        [7:0]    _zz_stateReg_31;
  reg        [7:0]    _zz_stateReg_32;
  reg        [7:0]    _zz_stateReg_33;
  reg        [7:0]    _zz_stateReg_34;
  reg        [7:0]    _zz_stateReg_35;
  wire                when_AES128_l192;
  wire       [7:0]    _zz_stateReg_36;
  wire       [7:0]    _zz_stateReg_37;
  wire       [7:0]    _zz_stateReg_38;
  wire       [7:0]    _zz_stateReg_39;
  wire       [7:0]    _zz_stateReg_40;
  wire       [7:0]    _zz_stateReg_41;
  wire       [7:0]    _zz_stateReg_42;
  wire       [7:0]    _zz_stateReg_43;
  wire       [7:0]    _zz_stateReg_44;
  wire       [7:0]    _zz_stateReg_45;
  wire       [7:0]    _zz_stateReg_46;
  wire       [7:0]    _zz_stateReg_47;
  wire       [7:0]    _zz_stateReg_48;
  wire       [7:0]    _zz_stateReg_49;
  wire       [7:0]    _zz_stateReg_50;
  wire       [7:0]    _zz_stateReg_51;
  wire       [7:0]    _zz_stateReg_52;
  wire       [7:0]    _zz_stateReg_53;
  wire       [7:0]    _zz_stateReg_54;
  wire       [7:0]    _zz_stateReg_55;
  wire       [7:0]    _zz_stateReg_56;
  wire       [7:0]    _zz_stateReg_57;
  wire       [7:0]    _zz_stateReg_58;
  wire       [7:0]    _zz_stateReg_59;
  wire       [7:0]    _zz_stateReg_60;
  wire       [7:0]    _zz_stateReg_61;
  wire       [7:0]    _zz_stateReg_62;
  wire       [7:0]    _zz_stateReg_63;
  wire       [7:0]    _zz_stateReg_64;
  wire       [7:0]    _zz_stateReg_65;
  wire       [7:0]    _zz_stateReg_66;
  wire       [7:0]    _zz_stateReg_67;
  wire       [127:0]  _zz_stateReg_68;
  wire       [31:0]   _zz_roundKeyReg_0;
  wire       [31:0]   _zz_roundKeyReg_0_1;
  wire       [31:0]   _zz_roundKeyReg_1;
  wire       [31:0]   _zz_roundKeyReg_2;
  wire       [31:0]   _zz_roundKeyReg_3;
  wire       [127:0]  _zz_stateReg_69;
  wire                when_AES128_l227;
  wire                when_AES128_l233;

  assign _zz__zz_stateReg_36 = ({1'd0,_zz_stateReg_4} <<< 1'd1);
  assign _zz__zz_stateReg_37 = ({1'd0,_zz_stateReg_5} <<< 1'd1);
  assign _zz__zz_stateReg_38 = ({1'd0,_zz_stateReg_5} <<< 1'd1);
  assign _zz__zz_stateReg_39 = ({1'd0,_zz_stateReg_6} <<< 1'd1);
  assign _zz__zz_stateReg_40 = ({1'd0,_zz_stateReg_6} <<< 1'd1);
  assign _zz__zz_stateReg_41 = ({1'd0,_zz_stateReg_7} <<< 1'd1);
  assign _zz__zz_stateReg_42 = ({1'd0,_zz_stateReg_4} <<< 1'd1);
  assign _zz__zz_stateReg_43 = ({1'd0,_zz_stateReg_7} <<< 1'd1);
  assign _zz__zz_stateReg_44 = ({1'd0,_zz_stateReg_8} <<< 1'd1);
  assign _zz__zz_stateReg_45 = ({1'd0,_zz_stateReg_9} <<< 1'd1);
  assign _zz__zz_stateReg_46 = ({1'd0,_zz_stateReg_9} <<< 1'd1);
  assign _zz__zz_stateReg_47 = ({1'd0,_zz_stateReg_10} <<< 1'd1);
  assign _zz__zz_stateReg_48 = ({1'd0,_zz_stateReg_10} <<< 1'd1);
  assign _zz__zz_stateReg_49 = ({1'd0,_zz_stateReg_11} <<< 1'd1);
  assign _zz__zz_stateReg_50 = ({1'd0,_zz_stateReg_8} <<< 1'd1);
  assign _zz__zz_stateReg_51 = ({1'd0,_zz_stateReg_11} <<< 1'd1);
  assign _zz__zz_stateReg_52 = ({1'd0,_zz_stateReg_12} <<< 1'd1);
  assign _zz__zz_stateReg_53 = ({1'd0,_zz_stateReg_13} <<< 1'd1);
  assign _zz__zz_stateReg_54 = ({1'd0,_zz_stateReg_13} <<< 1'd1);
  assign _zz__zz_stateReg_55 = ({1'd0,_zz_stateReg_14} <<< 1'd1);
  assign _zz__zz_stateReg_56 = ({1'd0,_zz_stateReg_14} <<< 1'd1);
  assign _zz__zz_stateReg_57 = ({1'd0,_zz_stateReg_15} <<< 1'd1);
  assign _zz__zz_stateReg_58 = ({1'd0,_zz_stateReg_12} <<< 1'd1);
  assign _zz__zz_stateReg_59 = ({1'd0,_zz_stateReg_15} <<< 1'd1);
  assign _zz__zz_stateReg_60 = ({1'd0,_zz_stateReg_16} <<< 1'd1);
  assign _zz__zz_stateReg_61 = ({1'd0,_zz_stateReg_17} <<< 1'd1);
  assign _zz__zz_stateReg_62 = ({1'd0,_zz_stateReg_17} <<< 1'd1);
  assign _zz__zz_stateReg_63 = ({1'd0,_zz_stateReg_18} <<< 1'd1);
  assign _zz__zz_stateReg_64 = ({1'd0,_zz_stateReg_18} <<< 1'd1);
  assign _zz__zz_stateReg_65 = ({1'd0,_zz_stateReg_19} <<< 1'd1);
  assign _zz__zz_stateReg_66 = ({1'd0,_zz_stateReg_16} <<< 1'd1);
  assign _zz__zz_stateReg_67 = ({1'd0,_zz_stateReg_19} <<< 1'd1);
  assign _zz__zz_stateReg_4_1 = stateReg[127 : 120];
  assign _zz__zz_stateReg_8_1 = stateReg[95 : 88];
  assign _zz__zz_stateReg_12_1 = stateReg[63 : 56];
  assign _zz__zz_stateReg_16_1 = stateReg[31 : 24];
  assign _zz__zz_stateReg_5_1 = stateReg[87 : 80];
  assign _zz__zz_stateReg_9_1 = stateReg[55 : 48];
  assign _zz__zz_stateReg_13_1 = stateReg[23 : 16];
  assign _zz__zz_stateReg_17_1 = stateReg[119 : 112];
  assign _zz__zz_stateReg_6_1 = stateReg[47 : 40];
  assign _zz__zz_stateReg_10_1 = stateReg[15 : 8];
  assign _zz__zz_stateReg_14_1 = stateReg[111 : 104];
  assign _zz__zz_stateReg_18_1 = stateReg[79 : 72];
  assign _zz__zz_stateReg_7_1 = stateReg[7 : 0];
  assign _zz__zz_stateReg_11_1 = stateReg[103 : 96];
  assign _zz__zz_stateReg_15_1 = stateReg[71 : 64];
  assign _zz__zz_stateReg_19_1 = stateReg[39 : 32];
  assign _zz__zz_roundKeyReg_0_1_1 = _zz_roundKeyReg_0[31 : 24];
  assign _zz__zz_roundKeyReg_0_1_3 = _zz_roundKeyReg_0[23 : 16];
  assign _zz__zz_roundKeyReg_0_1_5 = _zz_roundKeyReg_0[15 : 8];
  assign _zz__zz_roundKeyReg_0_1_7 = _zz_roundKeyReg_0[7 : 0];
  assign _zz_stateReg_70 = {{{{{_zz_stateReg_71,_zz_stateReg_77},_zz_stateReg_78},(_zz_stateReg_79 ^ _zz_stateReg_80)},(_zz_stateReg_81 ^ _zz_stateReg_2[31 : 24])},(io_dataIn[55 : 48] ^ _zz_stateReg_2[23 : 16])};
  assign _zz_stateReg_82 = (io_dataIn[47 : 40] ^ _zz_stateReg_2[15 : 8]);
  assign _zz_stateReg_83 = (io_dataIn[39 : 32] ^ _zz_stateReg_2[7 : 0]);
  assign _zz_stateReg_84 = io_dataIn[31 : 24];
  assign _zz_stateReg_85 = _zz_stateReg_3[31 : 24];
  assign _zz_stateReg_86 = io_dataIn[23 : 16];
  assign _zz_stateReg_71 = {{{{_zz_stateReg_72,_zz_stateReg_73},(_zz_stateReg_74 ^ _zz_stateReg_75)},(_zz_stateReg_76 ^ _zz_stateReg[7 : 0])},(io_dataIn[95 : 88] ^ _zz_stateReg_1[31 : 24])};
  assign _zz_stateReg_77 = (io_dataIn[87 : 80] ^ _zz_stateReg_1[23 : 16]);
  assign _zz_stateReg_78 = (io_dataIn[79 : 72] ^ _zz_stateReg_1[15 : 8]);
  assign _zz_stateReg_79 = io_dataIn[71 : 64];
  assign _zz_stateReg_80 = _zz_stateReg_1[7 : 0];
  assign _zz_stateReg_81 = io_dataIn[63 : 56];
  assign _zz_stateReg_72 = (io_dataIn[127 : 120] ^ _zz_stateReg[31 : 24]);
  assign _zz_stateReg_73 = (io_dataIn[119 : 112] ^ _zz_stateReg[23 : 16]);
  assign _zz_stateReg_74 = io_dataIn[111 : 104];
  assign _zz_stateReg_75 = _zz_stateReg[15 : 8];
  assign _zz_stateReg_76 = io_dataIn[103 : 96];
  assign _zz__zz_stateReg_68 = {{{{_zz_stateReg_20,_zz_stateReg_21},_zz_stateReg_22},_zz_stateReg_23},_zz_stateReg_24};
  assign _zz__zz_stateReg_68_1 = _zz_stateReg_25;
  assign _zz__zz_stateReg_69 = {{{{{{_zz_roundKeyReg_0_1[31 : 24],_zz_roundKeyReg_0_1[23 : 16]},_zz_roundKeyReg_0_1[15 : 8]},_zz_roundKeyReg_0_1[7 : 0]},_zz_roundKeyReg_1[31 : 24]},_zz_roundKeyReg_1[23 : 16]},_zz_roundKeyReg_1[15 : 8]};
  assign _zz__zz_stateReg_69_1 = _zz_roundKeyReg_1[7 : 0];
  assign _zz__zz_stateReg_69_2 = _zz_roundKeyReg_2[31 : 24];
  always @(*) begin
    case(_zz__zz_stateReg_4_1)
      8'b00000000 : _zz__zz_stateReg_4 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_4 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_4 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_4 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_4 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_4 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_4 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_4 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_4 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_4 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_4 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_4 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_4 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_4 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_4 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_4 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_4 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_4 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_4 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_4 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_4 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_4 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_4 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_4 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_4 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_4 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_4 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_4 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_4 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_4 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_4 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_4 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_4 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_4 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_4 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_4 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_4 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_4 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_4 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_4 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_4 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_4 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_4 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_4 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_4 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_4 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_4 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_4 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_4 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_4 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_4 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_4 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_4 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_4 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_4 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_4 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_4 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_4 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_4 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_4 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_4 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_4 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_4 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_4 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_4 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_4 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_4 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_4 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_4 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_4 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_4 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_4 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_4 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_4 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_4 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_4 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_4 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_4 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_4 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_4 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_4 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_4 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_4 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_4 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_4 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_4 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_4 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_4 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_4 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_4 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_4 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_4 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_4 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_4 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_4 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_4 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_4 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_4 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_4 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_4 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_4 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_4 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_4 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_4 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_4 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_4 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_4 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_4 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_4 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_4 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_4 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_4 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_4 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_4 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_4 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_4 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_4 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_4 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_4 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_4 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_4 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_4 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_4 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_4 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_4 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_4 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_4 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_4 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_4 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_4 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_4 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_4 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_4 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_4 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_4 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_4 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_4 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_4 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_4 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_4 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_4 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_4 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_4 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_4 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_4 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_4 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_4 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_4 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_4 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_4 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_4 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_4 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_4 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_4 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_4 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_4 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_4 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_4 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_4 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_4 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_4 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_4 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_4 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_4 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_4 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_4 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_4 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_4 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_4 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_4 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_4 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_4 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_4 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_4 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_4 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_4 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_4 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_4 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_4 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_4 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_4 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_4 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_4 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_4 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_4 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_4 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_4 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_4 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_4 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_4 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_4 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_4 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_4 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_4 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_4 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_4 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_4 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_4 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_4 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_4 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_4 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_4 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_4 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_4 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_4 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_4 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_4 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_4 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_4 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_4 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_4 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_4 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_4 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_4 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_4 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_4 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_4 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_4 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_4 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_4 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_4 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_4 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_4 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_4 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_4 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_4 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_4 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_4 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_4 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_4 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_4 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_4 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_4 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_4 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_4 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_4 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_4 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_4 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_4 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_4 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_4 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_4 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_4 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_4 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_4 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_4 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_4 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_4 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_4 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_4 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_4 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_4 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_4 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_4 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_4 = sboxRom_254;
      default : _zz__zz_stateReg_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_8_1)
      8'b00000000 : _zz__zz_stateReg_8 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_8 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_8 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_8 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_8 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_8 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_8 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_8 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_8 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_8 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_8 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_8 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_8 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_8 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_8 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_8 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_8 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_8 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_8 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_8 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_8 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_8 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_8 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_8 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_8 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_8 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_8 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_8 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_8 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_8 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_8 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_8 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_8 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_8 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_8 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_8 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_8 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_8 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_8 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_8 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_8 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_8 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_8 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_8 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_8 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_8 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_8 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_8 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_8 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_8 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_8 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_8 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_8 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_8 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_8 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_8 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_8 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_8 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_8 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_8 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_8 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_8 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_8 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_8 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_8 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_8 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_8 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_8 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_8 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_8 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_8 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_8 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_8 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_8 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_8 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_8 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_8 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_8 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_8 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_8 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_8 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_8 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_8 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_8 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_8 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_8 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_8 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_8 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_8 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_8 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_8 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_8 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_8 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_8 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_8 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_8 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_8 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_8 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_8 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_8 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_8 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_8 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_8 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_8 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_8 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_8 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_8 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_8 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_8 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_8 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_8 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_8 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_8 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_8 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_8 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_8 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_8 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_8 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_8 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_8 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_8 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_8 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_8 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_8 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_8 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_8 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_8 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_8 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_8 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_8 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_8 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_8 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_8 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_8 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_8 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_8 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_8 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_8 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_8 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_8 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_8 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_8 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_8 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_8 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_8 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_8 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_8 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_8 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_8 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_8 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_8 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_8 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_8 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_8 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_8 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_8 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_8 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_8 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_8 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_8 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_8 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_8 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_8 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_8 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_8 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_8 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_8 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_8 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_8 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_8 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_8 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_8 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_8 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_8 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_8 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_8 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_8 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_8 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_8 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_8 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_8 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_8 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_8 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_8 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_8 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_8 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_8 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_8 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_8 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_8 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_8 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_8 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_8 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_8 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_8 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_8 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_8 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_8 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_8 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_8 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_8 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_8 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_8 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_8 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_8 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_8 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_8 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_8 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_8 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_8 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_8 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_8 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_8 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_8 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_8 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_8 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_8 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_8 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_8 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_8 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_8 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_8 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_8 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_8 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_8 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_8 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_8 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_8 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_8 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_8 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_8 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_8 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_8 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_8 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_8 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_8 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_8 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_8 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_8 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_8 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_8 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_8 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_8 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_8 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_8 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_8 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_8 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_8 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_8 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_8 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_8 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_8 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_8 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_8 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_8 = sboxRom_254;
      default : _zz__zz_stateReg_8 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_12_1)
      8'b00000000 : _zz__zz_stateReg_12 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_12 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_12 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_12 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_12 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_12 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_12 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_12 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_12 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_12 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_12 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_12 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_12 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_12 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_12 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_12 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_12 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_12 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_12 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_12 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_12 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_12 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_12 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_12 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_12 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_12 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_12 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_12 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_12 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_12 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_12 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_12 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_12 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_12 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_12 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_12 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_12 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_12 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_12 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_12 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_12 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_12 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_12 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_12 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_12 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_12 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_12 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_12 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_12 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_12 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_12 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_12 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_12 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_12 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_12 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_12 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_12 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_12 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_12 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_12 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_12 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_12 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_12 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_12 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_12 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_12 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_12 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_12 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_12 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_12 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_12 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_12 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_12 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_12 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_12 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_12 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_12 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_12 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_12 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_12 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_12 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_12 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_12 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_12 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_12 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_12 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_12 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_12 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_12 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_12 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_12 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_12 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_12 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_12 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_12 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_12 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_12 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_12 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_12 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_12 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_12 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_12 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_12 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_12 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_12 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_12 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_12 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_12 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_12 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_12 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_12 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_12 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_12 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_12 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_12 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_12 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_12 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_12 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_12 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_12 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_12 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_12 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_12 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_12 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_12 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_12 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_12 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_12 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_12 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_12 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_12 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_12 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_12 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_12 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_12 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_12 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_12 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_12 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_12 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_12 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_12 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_12 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_12 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_12 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_12 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_12 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_12 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_12 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_12 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_12 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_12 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_12 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_12 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_12 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_12 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_12 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_12 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_12 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_12 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_12 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_12 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_12 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_12 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_12 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_12 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_12 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_12 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_12 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_12 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_12 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_12 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_12 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_12 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_12 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_12 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_12 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_12 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_12 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_12 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_12 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_12 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_12 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_12 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_12 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_12 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_12 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_12 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_12 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_12 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_12 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_12 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_12 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_12 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_12 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_12 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_12 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_12 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_12 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_12 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_12 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_12 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_12 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_12 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_12 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_12 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_12 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_12 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_12 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_12 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_12 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_12 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_12 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_12 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_12 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_12 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_12 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_12 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_12 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_12 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_12 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_12 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_12 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_12 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_12 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_12 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_12 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_12 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_12 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_12 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_12 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_12 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_12 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_12 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_12 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_12 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_12 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_12 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_12 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_12 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_12 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_12 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_12 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_12 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_12 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_12 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_12 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_12 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_12 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_12 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_12 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_12 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_12 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_12 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_12 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_12 = sboxRom_254;
      default : _zz__zz_stateReg_12 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_16_1)
      8'b00000000 : _zz__zz_stateReg_16 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_16 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_16 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_16 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_16 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_16 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_16 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_16 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_16 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_16 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_16 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_16 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_16 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_16 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_16 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_16 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_16 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_16 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_16 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_16 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_16 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_16 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_16 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_16 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_16 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_16 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_16 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_16 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_16 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_16 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_16 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_16 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_16 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_16 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_16 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_16 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_16 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_16 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_16 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_16 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_16 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_16 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_16 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_16 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_16 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_16 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_16 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_16 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_16 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_16 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_16 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_16 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_16 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_16 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_16 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_16 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_16 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_16 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_16 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_16 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_16 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_16 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_16 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_16 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_16 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_16 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_16 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_16 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_16 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_16 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_16 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_16 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_16 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_16 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_16 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_16 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_16 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_16 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_16 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_16 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_16 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_16 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_16 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_16 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_16 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_16 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_16 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_16 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_16 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_16 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_16 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_16 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_16 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_16 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_16 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_16 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_16 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_16 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_16 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_16 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_16 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_16 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_16 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_16 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_16 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_16 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_16 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_16 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_16 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_16 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_16 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_16 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_16 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_16 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_16 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_16 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_16 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_16 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_16 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_16 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_16 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_16 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_16 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_16 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_16 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_16 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_16 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_16 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_16 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_16 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_16 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_16 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_16 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_16 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_16 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_16 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_16 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_16 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_16 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_16 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_16 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_16 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_16 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_16 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_16 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_16 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_16 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_16 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_16 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_16 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_16 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_16 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_16 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_16 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_16 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_16 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_16 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_16 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_16 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_16 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_16 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_16 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_16 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_16 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_16 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_16 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_16 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_16 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_16 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_16 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_16 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_16 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_16 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_16 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_16 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_16 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_16 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_16 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_16 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_16 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_16 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_16 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_16 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_16 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_16 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_16 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_16 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_16 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_16 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_16 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_16 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_16 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_16 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_16 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_16 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_16 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_16 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_16 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_16 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_16 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_16 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_16 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_16 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_16 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_16 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_16 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_16 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_16 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_16 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_16 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_16 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_16 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_16 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_16 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_16 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_16 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_16 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_16 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_16 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_16 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_16 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_16 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_16 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_16 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_16 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_16 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_16 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_16 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_16 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_16 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_16 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_16 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_16 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_16 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_16 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_16 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_16 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_16 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_16 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_16 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_16 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_16 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_16 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_16 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_16 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_16 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_16 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_16 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_16 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_16 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_16 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_16 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_16 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_16 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_16 = sboxRom_254;
      default : _zz__zz_stateReg_16 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_5_1)
      8'b00000000 : _zz__zz_stateReg_5 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_5 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_5 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_5 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_5 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_5 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_5 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_5 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_5 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_5 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_5 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_5 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_5 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_5 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_5 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_5 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_5 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_5 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_5 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_5 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_5 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_5 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_5 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_5 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_5 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_5 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_5 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_5 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_5 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_5 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_5 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_5 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_5 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_5 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_5 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_5 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_5 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_5 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_5 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_5 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_5 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_5 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_5 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_5 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_5 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_5 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_5 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_5 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_5 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_5 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_5 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_5 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_5 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_5 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_5 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_5 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_5 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_5 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_5 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_5 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_5 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_5 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_5 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_5 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_5 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_5 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_5 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_5 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_5 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_5 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_5 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_5 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_5 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_5 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_5 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_5 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_5 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_5 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_5 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_5 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_5 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_5 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_5 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_5 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_5 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_5 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_5 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_5 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_5 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_5 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_5 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_5 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_5 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_5 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_5 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_5 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_5 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_5 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_5 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_5 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_5 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_5 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_5 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_5 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_5 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_5 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_5 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_5 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_5 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_5 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_5 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_5 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_5 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_5 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_5 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_5 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_5 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_5 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_5 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_5 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_5 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_5 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_5 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_5 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_5 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_5 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_5 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_5 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_5 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_5 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_5 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_5 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_5 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_5 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_5 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_5 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_5 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_5 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_5 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_5 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_5 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_5 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_5 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_5 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_5 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_5 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_5 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_5 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_5 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_5 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_5 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_5 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_5 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_5 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_5 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_5 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_5 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_5 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_5 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_5 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_5 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_5 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_5 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_5 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_5 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_5 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_5 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_5 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_5 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_5 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_5 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_5 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_5 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_5 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_5 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_5 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_5 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_5 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_5 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_5 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_5 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_5 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_5 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_5 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_5 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_5 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_5 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_5 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_5 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_5 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_5 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_5 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_5 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_5 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_5 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_5 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_5 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_5 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_5 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_5 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_5 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_5 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_5 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_5 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_5 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_5 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_5 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_5 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_5 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_5 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_5 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_5 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_5 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_5 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_5 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_5 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_5 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_5 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_5 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_5 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_5 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_5 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_5 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_5 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_5 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_5 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_5 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_5 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_5 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_5 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_5 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_5 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_5 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_5 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_5 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_5 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_5 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_5 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_5 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_5 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_5 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_5 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_5 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_5 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_5 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_5 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_5 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_5 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_5 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_5 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_5 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_5 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_5 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_5 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_5 = sboxRom_254;
      default : _zz__zz_stateReg_5 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_9_1)
      8'b00000000 : _zz__zz_stateReg_9 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_9 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_9 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_9 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_9 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_9 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_9 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_9 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_9 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_9 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_9 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_9 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_9 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_9 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_9 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_9 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_9 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_9 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_9 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_9 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_9 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_9 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_9 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_9 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_9 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_9 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_9 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_9 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_9 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_9 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_9 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_9 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_9 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_9 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_9 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_9 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_9 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_9 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_9 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_9 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_9 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_9 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_9 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_9 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_9 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_9 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_9 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_9 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_9 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_9 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_9 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_9 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_9 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_9 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_9 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_9 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_9 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_9 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_9 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_9 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_9 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_9 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_9 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_9 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_9 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_9 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_9 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_9 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_9 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_9 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_9 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_9 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_9 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_9 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_9 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_9 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_9 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_9 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_9 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_9 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_9 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_9 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_9 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_9 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_9 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_9 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_9 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_9 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_9 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_9 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_9 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_9 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_9 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_9 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_9 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_9 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_9 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_9 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_9 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_9 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_9 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_9 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_9 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_9 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_9 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_9 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_9 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_9 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_9 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_9 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_9 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_9 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_9 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_9 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_9 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_9 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_9 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_9 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_9 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_9 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_9 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_9 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_9 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_9 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_9 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_9 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_9 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_9 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_9 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_9 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_9 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_9 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_9 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_9 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_9 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_9 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_9 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_9 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_9 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_9 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_9 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_9 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_9 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_9 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_9 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_9 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_9 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_9 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_9 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_9 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_9 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_9 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_9 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_9 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_9 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_9 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_9 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_9 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_9 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_9 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_9 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_9 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_9 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_9 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_9 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_9 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_9 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_9 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_9 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_9 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_9 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_9 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_9 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_9 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_9 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_9 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_9 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_9 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_9 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_9 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_9 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_9 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_9 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_9 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_9 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_9 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_9 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_9 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_9 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_9 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_9 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_9 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_9 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_9 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_9 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_9 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_9 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_9 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_9 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_9 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_9 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_9 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_9 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_9 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_9 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_9 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_9 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_9 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_9 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_9 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_9 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_9 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_9 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_9 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_9 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_9 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_9 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_9 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_9 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_9 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_9 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_9 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_9 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_9 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_9 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_9 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_9 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_9 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_9 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_9 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_9 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_9 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_9 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_9 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_9 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_9 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_9 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_9 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_9 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_9 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_9 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_9 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_9 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_9 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_9 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_9 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_9 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_9 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_9 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_9 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_9 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_9 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_9 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_9 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_9 = sboxRom_254;
      default : _zz__zz_stateReg_9 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_13_1)
      8'b00000000 : _zz__zz_stateReg_13 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_13 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_13 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_13 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_13 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_13 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_13 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_13 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_13 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_13 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_13 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_13 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_13 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_13 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_13 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_13 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_13 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_13 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_13 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_13 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_13 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_13 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_13 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_13 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_13 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_13 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_13 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_13 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_13 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_13 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_13 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_13 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_13 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_13 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_13 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_13 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_13 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_13 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_13 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_13 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_13 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_13 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_13 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_13 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_13 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_13 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_13 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_13 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_13 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_13 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_13 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_13 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_13 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_13 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_13 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_13 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_13 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_13 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_13 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_13 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_13 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_13 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_13 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_13 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_13 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_13 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_13 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_13 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_13 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_13 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_13 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_13 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_13 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_13 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_13 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_13 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_13 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_13 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_13 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_13 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_13 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_13 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_13 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_13 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_13 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_13 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_13 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_13 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_13 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_13 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_13 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_13 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_13 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_13 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_13 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_13 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_13 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_13 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_13 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_13 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_13 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_13 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_13 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_13 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_13 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_13 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_13 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_13 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_13 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_13 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_13 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_13 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_13 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_13 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_13 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_13 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_13 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_13 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_13 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_13 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_13 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_13 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_13 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_13 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_13 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_13 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_13 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_13 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_13 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_13 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_13 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_13 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_13 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_13 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_13 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_13 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_13 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_13 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_13 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_13 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_13 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_13 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_13 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_13 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_13 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_13 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_13 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_13 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_13 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_13 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_13 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_13 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_13 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_13 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_13 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_13 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_13 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_13 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_13 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_13 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_13 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_13 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_13 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_13 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_13 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_13 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_13 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_13 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_13 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_13 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_13 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_13 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_13 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_13 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_13 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_13 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_13 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_13 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_13 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_13 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_13 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_13 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_13 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_13 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_13 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_13 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_13 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_13 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_13 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_13 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_13 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_13 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_13 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_13 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_13 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_13 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_13 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_13 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_13 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_13 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_13 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_13 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_13 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_13 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_13 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_13 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_13 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_13 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_13 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_13 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_13 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_13 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_13 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_13 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_13 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_13 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_13 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_13 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_13 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_13 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_13 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_13 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_13 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_13 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_13 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_13 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_13 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_13 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_13 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_13 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_13 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_13 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_13 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_13 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_13 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_13 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_13 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_13 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_13 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_13 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_13 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_13 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_13 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_13 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_13 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_13 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_13 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_13 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_13 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_13 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_13 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_13 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_13 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_13 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_13 = sboxRom_254;
      default : _zz__zz_stateReg_13 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_17_1)
      8'b00000000 : _zz__zz_stateReg_17 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_17 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_17 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_17 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_17 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_17 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_17 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_17 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_17 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_17 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_17 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_17 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_17 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_17 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_17 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_17 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_17 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_17 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_17 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_17 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_17 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_17 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_17 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_17 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_17 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_17 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_17 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_17 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_17 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_17 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_17 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_17 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_17 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_17 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_17 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_17 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_17 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_17 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_17 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_17 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_17 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_17 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_17 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_17 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_17 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_17 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_17 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_17 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_17 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_17 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_17 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_17 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_17 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_17 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_17 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_17 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_17 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_17 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_17 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_17 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_17 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_17 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_17 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_17 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_17 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_17 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_17 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_17 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_17 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_17 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_17 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_17 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_17 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_17 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_17 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_17 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_17 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_17 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_17 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_17 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_17 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_17 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_17 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_17 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_17 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_17 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_17 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_17 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_17 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_17 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_17 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_17 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_17 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_17 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_17 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_17 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_17 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_17 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_17 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_17 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_17 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_17 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_17 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_17 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_17 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_17 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_17 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_17 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_17 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_17 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_17 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_17 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_17 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_17 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_17 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_17 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_17 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_17 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_17 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_17 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_17 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_17 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_17 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_17 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_17 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_17 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_17 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_17 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_17 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_17 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_17 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_17 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_17 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_17 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_17 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_17 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_17 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_17 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_17 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_17 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_17 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_17 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_17 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_17 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_17 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_17 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_17 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_17 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_17 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_17 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_17 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_17 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_17 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_17 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_17 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_17 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_17 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_17 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_17 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_17 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_17 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_17 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_17 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_17 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_17 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_17 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_17 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_17 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_17 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_17 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_17 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_17 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_17 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_17 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_17 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_17 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_17 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_17 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_17 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_17 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_17 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_17 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_17 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_17 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_17 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_17 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_17 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_17 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_17 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_17 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_17 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_17 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_17 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_17 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_17 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_17 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_17 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_17 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_17 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_17 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_17 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_17 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_17 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_17 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_17 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_17 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_17 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_17 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_17 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_17 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_17 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_17 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_17 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_17 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_17 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_17 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_17 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_17 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_17 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_17 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_17 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_17 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_17 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_17 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_17 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_17 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_17 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_17 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_17 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_17 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_17 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_17 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_17 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_17 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_17 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_17 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_17 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_17 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_17 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_17 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_17 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_17 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_17 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_17 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_17 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_17 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_17 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_17 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_17 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_17 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_17 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_17 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_17 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_17 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_17 = sboxRom_254;
      default : _zz__zz_stateReg_17 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_6_1)
      8'b00000000 : _zz__zz_stateReg_6 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_6 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_6 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_6 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_6 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_6 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_6 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_6 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_6 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_6 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_6 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_6 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_6 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_6 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_6 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_6 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_6 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_6 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_6 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_6 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_6 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_6 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_6 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_6 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_6 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_6 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_6 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_6 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_6 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_6 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_6 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_6 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_6 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_6 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_6 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_6 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_6 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_6 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_6 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_6 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_6 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_6 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_6 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_6 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_6 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_6 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_6 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_6 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_6 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_6 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_6 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_6 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_6 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_6 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_6 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_6 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_6 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_6 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_6 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_6 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_6 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_6 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_6 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_6 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_6 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_6 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_6 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_6 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_6 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_6 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_6 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_6 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_6 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_6 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_6 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_6 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_6 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_6 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_6 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_6 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_6 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_6 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_6 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_6 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_6 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_6 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_6 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_6 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_6 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_6 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_6 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_6 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_6 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_6 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_6 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_6 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_6 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_6 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_6 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_6 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_6 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_6 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_6 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_6 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_6 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_6 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_6 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_6 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_6 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_6 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_6 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_6 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_6 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_6 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_6 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_6 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_6 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_6 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_6 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_6 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_6 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_6 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_6 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_6 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_6 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_6 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_6 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_6 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_6 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_6 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_6 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_6 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_6 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_6 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_6 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_6 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_6 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_6 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_6 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_6 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_6 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_6 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_6 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_6 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_6 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_6 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_6 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_6 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_6 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_6 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_6 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_6 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_6 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_6 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_6 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_6 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_6 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_6 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_6 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_6 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_6 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_6 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_6 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_6 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_6 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_6 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_6 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_6 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_6 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_6 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_6 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_6 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_6 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_6 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_6 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_6 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_6 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_6 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_6 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_6 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_6 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_6 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_6 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_6 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_6 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_6 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_6 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_6 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_6 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_6 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_6 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_6 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_6 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_6 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_6 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_6 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_6 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_6 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_6 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_6 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_6 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_6 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_6 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_6 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_6 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_6 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_6 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_6 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_6 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_6 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_6 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_6 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_6 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_6 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_6 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_6 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_6 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_6 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_6 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_6 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_6 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_6 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_6 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_6 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_6 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_6 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_6 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_6 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_6 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_6 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_6 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_6 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_6 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_6 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_6 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_6 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_6 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_6 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_6 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_6 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_6 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_6 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_6 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_6 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_6 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_6 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_6 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_6 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_6 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_6 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_6 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_6 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_6 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_6 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_6 = sboxRom_254;
      default : _zz__zz_stateReg_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_10_1)
      8'b00000000 : _zz__zz_stateReg_10 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_10 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_10 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_10 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_10 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_10 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_10 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_10 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_10 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_10 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_10 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_10 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_10 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_10 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_10 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_10 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_10 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_10 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_10 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_10 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_10 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_10 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_10 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_10 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_10 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_10 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_10 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_10 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_10 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_10 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_10 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_10 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_10 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_10 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_10 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_10 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_10 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_10 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_10 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_10 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_10 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_10 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_10 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_10 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_10 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_10 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_10 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_10 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_10 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_10 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_10 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_10 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_10 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_10 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_10 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_10 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_10 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_10 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_10 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_10 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_10 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_10 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_10 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_10 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_10 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_10 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_10 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_10 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_10 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_10 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_10 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_10 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_10 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_10 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_10 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_10 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_10 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_10 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_10 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_10 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_10 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_10 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_10 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_10 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_10 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_10 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_10 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_10 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_10 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_10 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_10 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_10 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_10 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_10 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_10 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_10 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_10 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_10 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_10 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_10 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_10 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_10 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_10 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_10 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_10 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_10 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_10 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_10 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_10 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_10 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_10 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_10 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_10 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_10 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_10 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_10 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_10 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_10 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_10 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_10 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_10 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_10 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_10 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_10 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_10 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_10 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_10 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_10 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_10 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_10 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_10 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_10 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_10 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_10 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_10 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_10 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_10 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_10 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_10 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_10 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_10 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_10 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_10 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_10 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_10 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_10 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_10 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_10 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_10 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_10 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_10 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_10 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_10 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_10 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_10 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_10 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_10 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_10 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_10 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_10 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_10 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_10 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_10 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_10 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_10 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_10 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_10 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_10 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_10 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_10 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_10 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_10 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_10 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_10 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_10 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_10 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_10 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_10 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_10 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_10 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_10 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_10 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_10 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_10 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_10 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_10 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_10 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_10 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_10 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_10 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_10 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_10 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_10 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_10 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_10 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_10 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_10 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_10 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_10 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_10 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_10 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_10 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_10 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_10 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_10 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_10 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_10 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_10 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_10 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_10 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_10 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_10 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_10 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_10 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_10 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_10 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_10 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_10 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_10 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_10 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_10 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_10 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_10 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_10 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_10 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_10 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_10 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_10 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_10 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_10 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_10 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_10 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_10 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_10 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_10 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_10 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_10 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_10 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_10 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_10 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_10 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_10 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_10 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_10 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_10 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_10 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_10 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_10 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_10 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_10 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_10 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_10 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_10 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_10 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_10 = sboxRom_254;
      default : _zz__zz_stateReg_10 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_14_1)
      8'b00000000 : _zz__zz_stateReg_14 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_14 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_14 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_14 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_14 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_14 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_14 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_14 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_14 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_14 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_14 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_14 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_14 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_14 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_14 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_14 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_14 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_14 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_14 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_14 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_14 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_14 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_14 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_14 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_14 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_14 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_14 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_14 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_14 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_14 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_14 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_14 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_14 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_14 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_14 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_14 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_14 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_14 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_14 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_14 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_14 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_14 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_14 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_14 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_14 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_14 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_14 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_14 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_14 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_14 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_14 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_14 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_14 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_14 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_14 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_14 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_14 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_14 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_14 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_14 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_14 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_14 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_14 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_14 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_14 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_14 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_14 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_14 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_14 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_14 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_14 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_14 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_14 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_14 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_14 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_14 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_14 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_14 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_14 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_14 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_14 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_14 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_14 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_14 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_14 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_14 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_14 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_14 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_14 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_14 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_14 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_14 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_14 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_14 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_14 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_14 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_14 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_14 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_14 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_14 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_14 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_14 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_14 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_14 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_14 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_14 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_14 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_14 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_14 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_14 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_14 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_14 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_14 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_14 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_14 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_14 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_14 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_14 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_14 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_14 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_14 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_14 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_14 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_14 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_14 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_14 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_14 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_14 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_14 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_14 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_14 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_14 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_14 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_14 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_14 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_14 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_14 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_14 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_14 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_14 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_14 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_14 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_14 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_14 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_14 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_14 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_14 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_14 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_14 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_14 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_14 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_14 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_14 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_14 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_14 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_14 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_14 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_14 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_14 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_14 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_14 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_14 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_14 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_14 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_14 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_14 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_14 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_14 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_14 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_14 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_14 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_14 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_14 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_14 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_14 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_14 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_14 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_14 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_14 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_14 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_14 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_14 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_14 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_14 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_14 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_14 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_14 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_14 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_14 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_14 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_14 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_14 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_14 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_14 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_14 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_14 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_14 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_14 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_14 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_14 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_14 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_14 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_14 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_14 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_14 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_14 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_14 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_14 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_14 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_14 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_14 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_14 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_14 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_14 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_14 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_14 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_14 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_14 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_14 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_14 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_14 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_14 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_14 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_14 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_14 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_14 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_14 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_14 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_14 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_14 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_14 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_14 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_14 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_14 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_14 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_14 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_14 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_14 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_14 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_14 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_14 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_14 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_14 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_14 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_14 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_14 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_14 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_14 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_14 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_14 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_14 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_14 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_14 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_14 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_14 = sboxRom_254;
      default : _zz__zz_stateReg_14 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_18_1)
      8'b00000000 : _zz__zz_stateReg_18 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_18 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_18 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_18 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_18 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_18 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_18 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_18 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_18 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_18 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_18 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_18 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_18 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_18 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_18 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_18 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_18 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_18 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_18 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_18 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_18 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_18 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_18 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_18 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_18 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_18 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_18 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_18 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_18 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_18 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_18 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_18 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_18 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_18 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_18 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_18 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_18 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_18 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_18 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_18 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_18 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_18 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_18 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_18 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_18 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_18 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_18 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_18 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_18 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_18 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_18 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_18 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_18 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_18 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_18 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_18 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_18 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_18 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_18 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_18 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_18 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_18 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_18 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_18 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_18 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_18 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_18 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_18 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_18 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_18 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_18 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_18 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_18 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_18 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_18 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_18 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_18 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_18 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_18 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_18 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_18 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_18 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_18 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_18 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_18 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_18 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_18 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_18 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_18 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_18 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_18 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_18 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_18 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_18 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_18 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_18 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_18 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_18 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_18 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_18 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_18 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_18 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_18 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_18 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_18 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_18 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_18 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_18 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_18 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_18 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_18 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_18 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_18 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_18 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_18 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_18 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_18 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_18 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_18 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_18 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_18 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_18 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_18 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_18 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_18 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_18 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_18 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_18 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_18 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_18 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_18 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_18 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_18 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_18 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_18 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_18 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_18 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_18 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_18 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_18 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_18 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_18 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_18 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_18 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_18 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_18 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_18 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_18 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_18 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_18 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_18 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_18 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_18 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_18 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_18 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_18 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_18 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_18 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_18 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_18 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_18 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_18 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_18 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_18 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_18 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_18 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_18 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_18 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_18 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_18 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_18 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_18 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_18 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_18 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_18 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_18 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_18 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_18 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_18 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_18 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_18 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_18 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_18 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_18 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_18 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_18 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_18 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_18 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_18 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_18 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_18 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_18 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_18 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_18 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_18 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_18 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_18 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_18 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_18 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_18 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_18 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_18 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_18 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_18 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_18 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_18 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_18 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_18 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_18 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_18 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_18 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_18 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_18 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_18 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_18 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_18 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_18 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_18 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_18 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_18 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_18 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_18 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_18 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_18 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_18 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_18 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_18 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_18 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_18 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_18 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_18 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_18 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_18 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_18 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_18 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_18 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_18 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_18 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_18 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_18 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_18 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_18 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_18 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_18 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_18 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_18 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_18 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_18 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_18 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_18 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_18 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_18 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_18 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_18 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_18 = sboxRom_254;
      default : _zz__zz_stateReg_18 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_7_1)
      8'b00000000 : _zz__zz_stateReg_7 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_7 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_7 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_7 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_7 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_7 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_7 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_7 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_7 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_7 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_7 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_7 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_7 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_7 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_7 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_7 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_7 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_7 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_7 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_7 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_7 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_7 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_7 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_7 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_7 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_7 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_7 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_7 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_7 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_7 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_7 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_7 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_7 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_7 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_7 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_7 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_7 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_7 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_7 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_7 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_7 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_7 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_7 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_7 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_7 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_7 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_7 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_7 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_7 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_7 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_7 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_7 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_7 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_7 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_7 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_7 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_7 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_7 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_7 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_7 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_7 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_7 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_7 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_7 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_7 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_7 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_7 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_7 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_7 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_7 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_7 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_7 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_7 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_7 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_7 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_7 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_7 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_7 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_7 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_7 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_7 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_7 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_7 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_7 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_7 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_7 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_7 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_7 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_7 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_7 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_7 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_7 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_7 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_7 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_7 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_7 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_7 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_7 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_7 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_7 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_7 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_7 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_7 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_7 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_7 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_7 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_7 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_7 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_7 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_7 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_7 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_7 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_7 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_7 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_7 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_7 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_7 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_7 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_7 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_7 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_7 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_7 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_7 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_7 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_7 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_7 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_7 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_7 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_7 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_7 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_7 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_7 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_7 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_7 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_7 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_7 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_7 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_7 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_7 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_7 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_7 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_7 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_7 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_7 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_7 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_7 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_7 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_7 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_7 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_7 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_7 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_7 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_7 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_7 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_7 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_7 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_7 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_7 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_7 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_7 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_7 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_7 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_7 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_7 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_7 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_7 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_7 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_7 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_7 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_7 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_7 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_7 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_7 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_7 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_7 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_7 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_7 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_7 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_7 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_7 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_7 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_7 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_7 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_7 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_7 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_7 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_7 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_7 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_7 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_7 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_7 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_7 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_7 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_7 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_7 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_7 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_7 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_7 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_7 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_7 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_7 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_7 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_7 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_7 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_7 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_7 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_7 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_7 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_7 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_7 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_7 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_7 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_7 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_7 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_7 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_7 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_7 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_7 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_7 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_7 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_7 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_7 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_7 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_7 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_7 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_7 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_7 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_7 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_7 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_7 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_7 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_7 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_7 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_7 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_7 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_7 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_7 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_7 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_7 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_7 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_7 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_7 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_7 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_7 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_7 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_7 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_7 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_7 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_7 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_7 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_7 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_7 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_7 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_7 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_7 = sboxRom_254;
      default : _zz__zz_stateReg_7 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_11_1)
      8'b00000000 : _zz__zz_stateReg_11 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_11 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_11 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_11 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_11 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_11 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_11 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_11 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_11 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_11 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_11 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_11 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_11 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_11 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_11 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_11 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_11 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_11 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_11 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_11 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_11 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_11 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_11 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_11 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_11 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_11 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_11 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_11 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_11 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_11 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_11 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_11 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_11 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_11 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_11 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_11 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_11 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_11 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_11 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_11 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_11 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_11 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_11 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_11 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_11 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_11 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_11 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_11 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_11 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_11 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_11 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_11 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_11 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_11 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_11 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_11 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_11 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_11 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_11 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_11 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_11 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_11 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_11 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_11 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_11 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_11 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_11 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_11 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_11 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_11 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_11 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_11 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_11 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_11 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_11 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_11 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_11 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_11 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_11 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_11 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_11 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_11 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_11 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_11 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_11 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_11 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_11 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_11 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_11 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_11 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_11 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_11 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_11 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_11 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_11 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_11 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_11 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_11 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_11 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_11 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_11 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_11 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_11 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_11 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_11 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_11 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_11 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_11 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_11 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_11 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_11 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_11 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_11 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_11 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_11 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_11 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_11 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_11 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_11 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_11 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_11 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_11 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_11 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_11 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_11 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_11 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_11 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_11 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_11 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_11 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_11 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_11 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_11 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_11 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_11 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_11 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_11 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_11 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_11 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_11 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_11 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_11 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_11 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_11 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_11 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_11 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_11 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_11 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_11 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_11 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_11 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_11 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_11 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_11 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_11 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_11 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_11 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_11 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_11 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_11 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_11 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_11 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_11 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_11 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_11 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_11 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_11 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_11 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_11 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_11 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_11 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_11 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_11 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_11 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_11 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_11 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_11 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_11 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_11 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_11 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_11 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_11 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_11 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_11 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_11 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_11 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_11 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_11 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_11 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_11 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_11 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_11 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_11 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_11 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_11 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_11 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_11 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_11 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_11 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_11 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_11 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_11 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_11 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_11 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_11 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_11 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_11 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_11 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_11 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_11 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_11 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_11 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_11 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_11 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_11 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_11 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_11 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_11 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_11 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_11 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_11 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_11 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_11 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_11 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_11 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_11 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_11 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_11 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_11 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_11 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_11 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_11 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_11 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_11 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_11 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_11 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_11 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_11 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_11 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_11 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_11 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_11 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_11 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_11 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_11 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_11 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_11 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_11 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_11 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_11 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_11 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_11 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_11 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_11 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_11 = sboxRom_254;
      default : _zz__zz_stateReg_11 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_15_1)
      8'b00000000 : _zz__zz_stateReg_15 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_15 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_15 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_15 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_15 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_15 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_15 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_15 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_15 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_15 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_15 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_15 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_15 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_15 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_15 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_15 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_15 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_15 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_15 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_15 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_15 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_15 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_15 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_15 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_15 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_15 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_15 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_15 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_15 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_15 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_15 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_15 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_15 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_15 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_15 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_15 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_15 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_15 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_15 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_15 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_15 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_15 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_15 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_15 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_15 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_15 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_15 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_15 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_15 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_15 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_15 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_15 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_15 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_15 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_15 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_15 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_15 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_15 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_15 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_15 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_15 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_15 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_15 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_15 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_15 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_15 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_15 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_15 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_15 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_15 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_15 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_15 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_15 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_15 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_15 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_15 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_15 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_15 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_15 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_15 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_15 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_15 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_15 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_15 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_15 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_15 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_15 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_15 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_15 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_15 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_15 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_15 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_15 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_15 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_15 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_15 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_15 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_15 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_15 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_15 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_15 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_15 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_15 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_15 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_15 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_15 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_15 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_15 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_15 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_15 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_15 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_15 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_15 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_15 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_15 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_15 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_15 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_15 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_15 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_15 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_15 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_15 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_15 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_15 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_15 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_15 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_15 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_15 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_15 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_15 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_15 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_15 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_15 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_15 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_15 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_15 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_15 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_15 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_15 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_15 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_15 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_15 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_15 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_15 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_15 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_15 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_15 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_15 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_15 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_15 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_15 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_15 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_15 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_15 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_15 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_15 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_15 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_15 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_15 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_15 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_15 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_15 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_15 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_15 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_15 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_15 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_15 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_15 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_15 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_15 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_15 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_15 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_15 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_15 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_15 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_15 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_15 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_15 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_15 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_15 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_15 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_15 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_15 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_15 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_15 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_15 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_15 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_15 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_15 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_15 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_15 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_15 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_15 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_15 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_15 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_15 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_15 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_15 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_15 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_15 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_15 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_15 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_15 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_15 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_15 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_15 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_15 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_15 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_15 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_15 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_15 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_15 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_15 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_15 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_15 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_15 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_15 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_15 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_15 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_15 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_15 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_15 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_15 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_15 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_15 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_15 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_15 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_15 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_15 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_15 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_15 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_15 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_15 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_15 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_15 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_15 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_15 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_15 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_15 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_15 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_15 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_15 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_15 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_15 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_15 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_15 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_15 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_15 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_15 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_15 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_15 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_15 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_15 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_15 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_15 = sboxRom_254;
      default : _zz__zz_stateReg_15 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_stateReg_19_1)
      8'b00000000 : _zz__zz_stateReg_19 = sboxRom_0;
      8'b00000001 : _zz__zz_stateReg_19 = sboxRom_1;
      8'b00000010 : _zz__zz_stateReg_19 = sboxRom_2;
      8'b00000011 : _zz__zz_stateReg_19 = sboxRom_3;
      8'b00000100 : _zz__zz_stateReg_19 = sboxRom_4;
      8'b00000101 : _zz__zz_stateReg_19 = sboxRom_5;
      8'b00000110 : _zz__zz_stateReg_19 = sboxRom_6;
      8'b00000111 : _zz__zz_stateReg_19 = sboxRom_7;
      8'b00001000 : _zz__zz_stateReg_19 = sboxRom_8;
      8'b00001001 : _zz__zz_stateReg_19 = sboxRom_9;
      8'b00001010 : _zz__zz_stateReg_19 = sboxRom_10;
      8'b00001011 : _zz__zz_stateReg_19 = sboxRom_11;
      8'b00001100 : _zz__zz_stateReg_19 = sboxRom_12;
      8'b00001101 : _zz__zz_stateReg_19 = sboxRom_13;
      8'b00001110 : _zz__zz_stateReg_19 = sboxRom_14;
      8'b00001111 : _zz__zz_stateReg_19 = sboxRom_15;
      8'b00010000 : _zz__zz_stateReg_19 = sboxRom_16;
      8'b00010001 : _zz__zz_stateReg_19 = sboxRom_17;
      8'b00010010 : _zz__zz_stateReg_19 = sboxRom_18;
      8'b00010011 : _zz__zz_stateReg_19 = sboxRom_19;
      8'b00010100 : _zz__zz_stateReg_19 = sboxRom_20;
      8'b00010101 : _zz__zz_stateReg_19 = sboxRom_21;
      8'b00010110 : _zz__zz_stateReg_19 = sboxRom_22;
      8'b00010111 : _zz__zz_stateReg_19 = sboxRom_23;
      8'b00011000 : _zz__zz_stateReg_19 = sboxRom_24;
      8'b00011001 : _zz__zz_stateReg_19 = sboxRom_25;
      8'b00011010 : _zz__zz_stateReg_19 = sboxRom_26;
      8'b00011011 : _zz__zz_stateReg_19 = sboxRom_27;
      8'b00011100 : _zz__zz_stateReg_19 = sboxRom_28;
      8'b00011101 : _zz__zz_stateReg_19 = sboxRom_29;
      8'b00011110 : _zz__zz_stateReg_19 = sboxRom_30;
      8'b00011111 : _zz__zz_stateReg_19 = sboxRom_31;
      8'b00100000 : _zz__zz_stateReg_19 = sboxRom_32;
      8'b00100001 : _zz__zz_stateReg_19 = sboxRom_33;
      8'b00100010 : _zz__zz_stateReg_19 = sboxRom_34;
      8'b00100011 : _zz__zz_stateReg_19 = sboxRom_35;
      8'b00100100 : _zz__zz_stateReg_19 = sboxRom_36;
      8'b00100101 : _zz__zz_stateReg_19 = sboxRom_37;
      8'b00100110 : _zz__zz_stateReg_19 = sboxRom_38;
      8'b00100111 : _zz__zz_stateReg_19 = sboxRom_39;
      8'b00101000 : _zz__zz_stateReg_19 = sboxRom_40;
      8'b00101001 : _zz__zz_stateReg_19 = sboxRom_41;
      8'b00101010 : _zz__zz_stateReg_19 = sboxRom_42;
      8'b00101011 : _zz__zz_stateReg_19 = sboxRom_43;
      8'b00101100 : _zz__zz_stateReg_19 = sboxRom_44;
      8'b00101101 : _zz__zz_stateReg_19 = sboxRom_45;
      8'b00101110 : _zz__zz_stateReg_19 = sboxRom_46;
      8'b00101111 : _zz__zz_stateReg_19 = sboxRom_47;
      8'b00110000 : _zz__zz_stateReg_19 = sboxRom_48;
      8'b00110001 : _zz__zz_stateReg_19 = sboxRom_49;
      8'b00110010 : _zz__zz_stateReg_19 = sboxRom_50;
      8'b00110011 : _zz__zz_stateReg_19 = sboxRom_51;
      8'b00110100 : _zz__zz_stateReg_19 = sboxRom_52;
      8'b00110101 : _zz__zz_stateReg_19 = sboxRom_53;
      8'b00110110 : _zz__zz_stateReg_19 = sboxRom_54;
      8'b00110111 : _zz__zz_stateReg_19 = sboxRom_55;
      8'b00111000 : _zz__zz_stateReg_19 = sboxRom_56;
      8'b00111001 : _zz__zz_stateReg_19 = sboxRom_57;
      8'b00111010 : _zz__zz_stateReg_19 = sboxRom_58;
      8'b00111011 : _zz__zz_stateReg_19 = sboxRom_59;
      8'b00111100 : _zz__zz_stateReg_19 = sboxRom_60;
      8'b00111101 : _zz__zz_stateReg_19 = sboxRom_61;
      8'b00111110 : _zz__zz_stateReg_19 = sboxRom_62;
      8'b00111111 : _zz__zz_stateReg_19 = sboxRom_63;
      8'b01000000 : _zz__zz_stateReg_19 = sboxRom_64;
      8'b01000001 : _zz__zz_stateReg_19 = sboxRom_65;
      8'b01000010 : _zz__zz_stateReg_19 = sboxRom_66;
      8'b01000011 : _zz__zz_stateReg_19 = sboxRom_67;
      8'b01000100 : _zz__zz_stateReg_19 = sboxRom_68;
      8'b01000101 : _zz__zz_stateReg_19 = sboxRom_69;
      8'b01000110 : _zz__zz_stateReg_19 = sboxRom_70;
      8'b01000111 : _zz__zz_stateReg_19 = sboxRom_71;
      8'b01001000 : _zz__zz_stateReg_19 = sboxRom_72;
      8'b01001001 : _zz__zz_stateReg_19 = sboxRom_73;
      8'b01001010 : _zz__zz_stateReg_19 = sboxRom_74;
      8'b01001011 : _zz__zz_stateReg_19 = sboxRom_75;
      8'b01001100 : _zz__zz_stateReg_19 = sboxRom_76;
      8'b01001101 : _zz__zz_stateReg_19 = sboxRom_77;
      8'b01001110 : _zz__zz_stateReg_19 = sboxRom_78;
      8'b01001111 : _zz__zz_stateReg_19 = sboxRom_79;
      8'b01010000 : _zz__zz_stateReg_19 = sboxRom_80;
      8'b01010001 : _zz__zz_stateReg_19 = sboxRom_81;
      8'b01010010 : _zz__zz_stateReg_19 = sboxRom_82;
      8'b01010011 : _zz__zz_stateReg_19 = sboxRom_83;
      8'b01010100 : _zz__zz_stateReg_19 = sboxRom_84;
      8'b01010101 : _zz__zz_stateReg_19 = sboxRom_85;
      8'b01010110 : _zz__zz_stateReg_19 = sboxRom_86;
      8'b01010111 : _zz__zz_stateReg_19 = sboxRom_87;
      8'b01011000 : _zz__zz_stateReg_19 = sboxRom_88;
      8'b01011001 : _zz__zz_stateReg_19 = sboxRom_89;
      8'b01011010 : _zz__zz_stateReg_19 = sboxRom_90;
      8'b01011011 : _zz__zz_stateReg_19 = sboxRom_91;
      8'b01011100 : _zz__zz_stateReg_19 = sboxRom_92;
      8'b01011101 : _zz__zz_stateReg_19 = sboxRom_93;
      8'b01011110 : _zz__zz_stateReg_19 = sboxRom_94;
      8'b01011111 : _zz__zz_stateReg_19 = sboxRom_95;
      8'b01100000 : _zz__zz_stateReg_19 = sboxRom_96;
      8'b01100001 : _zz__zz_stateReg_19 = sboxRom_97;
      8'b01100010 : _zz__zz_stateReg_19 = sboxRom_98;
      8'b01100011 : _zz__zz_stateReg_19 = sboxRom_99;
      8'b01100100 : _zz__zz_stateReg_19 = sboxRom_100;
      8'b01100101 : _zz__zz_stateReg_19 = sboxRom_101;
      8'b01100110 : _zz__zz_stateReg_19 = sboxRom_102;
      8'b01100111 : _zz__zz_stateReg_19 = sboxRom_103;
      8'b01101000 : _zz__zz_stateReg_19 = sboxRom_104;
      8'b01101001 : _zz__zz_stateReg_19 = sboxRom_105;
      8'b01101010 : _zz__zz_stateReg_19 = sboxRom_106;
      8'b01101011 : _zz__zz_stateReg_19 = sboxRom_107;
      8'b01101100 : _zz__zz_stateReg_19 = sboxRom_108;
      8'b01101101 : _zz__zz_stateReg_19 = sboxRom_109;
      8'b01101110 : _zz__zz_stateReg_19 = sboxRom_110;
      8'b01101111 : _zz__zz_stateReg_19 = sboxRom_111;
      8'b01110000 : _zz__zz_stateReg_19 = sboxRom_112;
      8'b01110001 : _zz__zz_stateReg_19 = sboxRom_113;
      8'b01110010 : _zz__zz_stateReg_19 = sboxRom_114;
      8'b01110011 : _zz__zz_stateReg_19 = sboxRom_115;
      8'b01110100 : _zz__zz_stateReg_19 = sboxRom_116;
      8'b01110101 : _zz__zz_stateReg_19 = sboxRom_117;
      8'b01110110 : _zz__zz_stateReg_19 = sboxRom_118;
      8'b01110111 : _zz__zz_stateReg_19 = sboxRom_119;
      8'b01111000 : _zz__zz_stateReg_19 = sboxRom_120;
      8'b01111001 : _zz__zz_stateReg_19 = sboxRom_121;
      8'b01111010 : _zz__zz_stateReg_19 = sboxRom_122;
      8'b01111011 : _zz__zz_stateReg_19 = sboxRom_123;
      8'b01111100 : _zz__zz_stateReg_19 = sboxRom_124;
      8'b01111101 : _zz__zz_stateReg_19 = sboxRom_125;
      8'b01111110 : _zz__zz_stateReg_19 = sboxRom_126;
      8'b01111111 : _zz__zz_stateReg_19 = sboxRom_127;
      8'b10000000 : _zz__zz_stateReg_19 = sboxRom_128;
      8'b10000001 : _zz__zz_stateReg_19 = sboxRom_129;
      8'b10000010 : _zz__zz_stateReg_19 = sboxRom_130;
      8'b10000011 : _zz__zz_stateReg_19 = sboxRom_131;
      8'b10000100 : _zz__zz_stateReg_19 = sboxRom_132;
      8'b10000101 : _zz__zz_stateReg_19 = sboxRom_133;
      8'b10000110 : _zz__zz_stateReg_19 = sboxRom_134;
      8'b10000111 : _zz__zz_stateReg_19 = sboxRom_135;
      8'b10001000 : _zz__zz_stateReg_19 = sboxRom_136;
      8'b10001001 : _zz__zz_stateReg_19 = sboxRom_137;
      8'b10001010 : _zz__zz_stateReg_19 = sboxRom_138;
      8'b10001011 : _zz__zz_stateReg_19 = sboxRom_139;
      8'b10001100 : _zz__zz_stateReg_19 = sboxRom_140;
      8'b10001101 : _zz__zz_stateReg_19 = sboxRom_141;
      8'b10001110 : _zz__zz_stateReg_19 = sboxRom_142;
      8'b10001111 : _zz__zz_stateReg_19 = sboxRom_143;
      8'b10010000 : _zz__zz_stateReg_19 = sboxRom_144;
      8'b10010001 : _zz__zz_stateReg_19 = sboxRom_145;
      8'b10010010 : _zz__zz_stateReg_19 = sboxRom_146;
      8'b10010011 : _zz__zz_stateReg_19 = sboxRom_147;
      8'b10010100 : _zz__zz_stateReg_19 = sboxRom_148;
      8'b10010101 : _zz__zz_stateReg_19 = sboxRom_149;
      8'b10010110 : _zz__zz_stateReg_19 = sboxRom_150;
      8'b10010111 : _zz__zz_stateReg_19 = sboxRom_151;
      8'b10011000 : _zz__zz_stateReg_19 = sboxRom_152;
      8'b10011001 : _zz__zz_stateReg_19 = sboxRom_153;
      8'b10011010 : _zz__zz_stateReg_19 = sboxRom_154;
      8'b10011011 : _zz__zz_stateReg_19 = sboxRom_155;
      8'b10011100 : _zz__zz_stateReg_19 = sboxRom_156;
      8'b10011101 : _zz__zz_stateReg_19 = sboxRom_157;
      8'b10011110 : _zz__zz_stateReg_19 = sboxRom_158;
      8'b10011111 : _zz__zz_stateReg_19 = sboxRom_159;
      8'b10100000 : _zz__zz_stateReg_19 = sboxRom_160;
      8'b10100001 : _zz__zz_stateReg_19 = sboxRom_161;
      8'b10100010 : _zz__zz_stateReg_19 = sboxRom_162;
      8'b10100011 : _zz__zz_stateReg_19 = sboxRom_163;
      8'b10100100 : _zz__zz_stateReg_19 = sboxRom_164;
      8'b10100101 : _zz__zz_stateReg_19 = sboxRom_165;
      8'b10100110 : _zz__zz_stateReg_19 = sboxRom_166;
      8'b10100111 : _zz__zz_stateReg_19 = sboxRom_167;
      8'b10101000 : _zz__zz_stateReg_19 = sboxRom_168;
      8'b10101001 : _zz__zz_stateReg_19 = sboxRom_169;
      8'b10101010 : _zz__zz_stateReg_19 = sboxRom_170;
      8'b10101011 : _zz__zz_stateReg_19 = sboxRom_171;
      8'b10101100 : _zz__zz_stateReg_19 = sboxRom_172;
      8'b10101101 : _zz__zz_stateReg_19 = sboxRom_173;
      8'b10101110 : _zz__zz_stateReg_19 = sboxRom_174;
      8'b10101111 : _zz__zz_stateReg_19 = sboxRom_175;
      8'b10110000 : _zz__zz_stateReg_19 = sboxRom_176;
      8'b10110001 : _zz__zz_stateReg_19 = sboxRom_177;
      8'b10110010 : _zz__zz_stateReg_19 = sboxRom_178;
      8'b10110011 : _zz__zz_stateReg_19 = sboxRom_179;
      8'b10110100 : _zz__zz_stateReg_19 = sboxRom_180;
      8'b10110101 : _zz__zz_stateReg_19 = sboxRom_181;
      8'b10110110 : _zz__zz_stateReg_19 = sboxRom_182;
      8'b10110111 : _zz__zz_stateReg_19 = sboxRom_183;
      8'b10111000 : _zz__zz_stateReg_19 = sboxRom_184;
      8'b10111001 : _zz__zz_stateReg_19 = sboxRom_185;
      8'b10111010 : _zz__zz_stateReg_19 = sboxRom_186;
      8'b10111011 : _zz__zz_stateReg_19 = sboxRom_187;
      8'b10111100 : _zz__zz_stateReg_19 = sboxRom_188;
      8'b10111101 : _zz__zz_stateReg_19 = sboxRom_189;
      8'b10111110 : _zz__zz_stateReg_19 = sboxRom_190;
      8'b10111111 : _zz__zz_stateReg_19 = sboxRom_191;
      8'b11000000 : _zz__zz_stateReg_19 = sboxRom_192;
      8'b11000001 : _zz__zz_stateReg_19 = sboxRom_193;
      8'b11000010 : _zz__zz_stateReg_19 = sboxRom_194;
      8'b11000011 : _zz__zz_stateReg_19 = sboxRom_195;
      8'b11000100 : _zz__zz_stateReg_19 = sboxRom_196;
      8'b11000101 : _zz__zz_stateReg_19 = sboxRom_197;
      8'b11000110 : _zz__zz_stateReg_19 = sboxRom_198;
      8'b11000111 : _zz__zz_stateReg_19 = sboxRom_199;
      8'b11001000 : _zz__zz_stateReg_19 = sboxRom_200;
      8'b11001001 : _zz__zz_stateReg_19 = sboxRom_201;
      8'b11001010 : _zz__zz_stateReg_19 = sboxRom_202;
      8'b11001011 : _zz__zz_stateReg_19 = sboxRom_203;
      8'b11001100 : _zz__zz_stateReg_19 = sboxRom_204;
      8'b11001101 : _zz__zz_stateReg_19 = sboxRom_205;
      8'b11001110 : _zz__zz_stateReg_19 = sboxRom_206;
      8'b11001111 : _zz__zz_stateReg_19 = sboxRom_207;
      8'b11010000 : _zz__zz_stateReg_19 = sboxRom_208;
      8'b11010001 : _zz__zz_stateReg_19 = sboxRom_209;
      8'b11010010 : _zz__zz_stateReg_19 = sboxRom_210;
      8'b11010011 : _zz__zz_stateReg_19 = sboxRom_211;
      8'b11010100 : _zz__zz_stateReg_19 = sboxRom_212;
      8'b11010101 : _zz__zz_stateReg_19 = sboxRom_213;
      8'b11010110 : _zz__zz_stateReg_19 = sboxRom_214;
      8'b11010111 : _zz__zz_stateReg_19 = sboxRom_215;
      8'b11011000 : _zz__zz_stateReg_19 = sboxRom_216;
      8'b11011001 : _zz__zz_stateReg_19 = sboxRom_217;
      8'b11011010 : _zz__zz_stateReg_19 = sboxRom_218;
      8'b11011011 : _zz__zz_stateReg_19 = sboxRom_219;
      8'b11011100 : _zz__zz_stateReg_19 = sboxRom_220;
      8'b11011101 : _zz__zz_stateReg_19 = sboxRom_221;
      8'b11011110 : _zz__zz_stateReg_19 = sboxRom_222;
      8'b11011111 : _zz__zz_stateReg_19 = sboxRom_223;
      8'b11100000 : _zz__zz_stateReg_19 = sboxRom_224;
      8'b11100001 : _zz__zz_stateReg_19 = sboxRom_225;
      8'b11100010 : _zz__zz_stateReg_19 = sboxRom_226;
      8'b11100011 : _zz__zz_stateReg_19 = sboxRom_227;
      8'b11100100 : _zz__zz_stateReg_19 = sboxRom_228;
      8'b11100101 : _zz__zz_stateReg_19 = sboxRom_229;
      8'b11100110 : _zz__zz_stateReg_19 = sboxRom_230;
      8'b11100111 : _zz__zz_stateReg_19 = sboxRom_231;
      8'b11101000 : _zz__zz_stateReg_19 = sboxRom_232;
      8'b11101001 : _zz__zz_stateReg_19 = sboxRom_233;
      8'b11101010 : _zz__zz_stateReg_19 = sboxRom_234;
      8'b11101011 : _zz__zz_stateReg_19 = sboxRom_235;
      8'b11101100 : _zz__zz_stateReg_19 = sboxRom_236;
      8'b11101101 : _zz__zz_stateReg_19 = sboxRom_237;
      8'b11101110 : _zz__zz_stateReg_19 = sboxRom_238;
      8'b11101111 : _zz__zz_stateReg_19 = sboxRom_239;
      8'b11110000 : _zz__zz_stateReg_19 = sboxRom_240;
      8'b11110001 : _zz__zz_stateReg_19 = sboxRom_241;
      8'b11110010 : _zz__zz_stateReg_19 = sboxRom_242;
      8'b11110011 : _zz__zz_stateReg_19 = sboxRom_243;
      8'b11110100 : _zz__zz_stateReg_19 = sboxRom_244;
      8'b11110101 : _zz__zz_stateReg_19 = sboxRom_245;
      8'b11110110 : _zz__zz_stateReg_19 = sboxRom_246;
      8'b11110111 : _zz__zz_stateReg_19 = sboxRom_247;
      8'b11111000 : _zz__zz_stateReg_19 = sboxRom_248;
      8'b11111001 : _zz__zz_stateReg_19 = sboxRom_249;
      8'b11111010 : _zz__zz_stateReg_19 = sboxRom_250;
      8'b11111011 : _zz__zz_stateReg_19 = sboxRom_251;
      8'b11111100 : _zz__zz_stateReg_19 = sboxRom_252;
      8'b11111101 : _zz__zz_stateReg_19 = sboxRom_253;
      8'b11111110 : _zz__zz_stateReg_19 = sboxRom_254;
      default : _zz__zz_stateReg_19 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_1_1)
      8'b00000000 : _zz__zz_roundKeyReg_0_1 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_1 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_1 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_1 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_1 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_1 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_1 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_1 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_1 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_1 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_1 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_1 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_1 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_1 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_1 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_1 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_1 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_1 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_1 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_1 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_1 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_1 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_1 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_1 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_1 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_1 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_1 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_1 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_1 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_1 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_1 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_1 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_1 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_1 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_1 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_1 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_1 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_1 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_1 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_1 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_1 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_1 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_1 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_1 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_1 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_1 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_1 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_1 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_1 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_1 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_1 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_1 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_1 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_1 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_1 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_1 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_1 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_1 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_1 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_1 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_1 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_1 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_1 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_1 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_1 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_1 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_1 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_1 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_1 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_1 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_1 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_1 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_1 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_1 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_1 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_1 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_1 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_1 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_1 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_1 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_1 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_1 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_1 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_1 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_1 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_1 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_1 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_1 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_1 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_1 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_1 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_1 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_1 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_1 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_1 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_1 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_1 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_1 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_1 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_1 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_1 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_1 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_1 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_1 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_1 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_1 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_1 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_1 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_1 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_1 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_1 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_1 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_1 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_1 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_1 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_1 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_1 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_1 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_1 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_1 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_1 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_1 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_1 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_1 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_1 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_1 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_1 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_1 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_1 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_1 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_1 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_1 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_1 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_1 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_1 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_1 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_1 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_1 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_1 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_1 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_1 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_1 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_1 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_1 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_1 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_1 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_1 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_1 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_1 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_1 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_1 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_1 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_1 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_1 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_1 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_1 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_1 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_1 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_1 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_1 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_1 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_1 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_1 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_1 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_1 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_1 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_1 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_1 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_1 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_1 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_1 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_1 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_1 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_1 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_1 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_1 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_1 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_1 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_1 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_1 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_1 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_1 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_1 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_1 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_1 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_1 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_1 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_1 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_1 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_1 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_1 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_1 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_1 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_1 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_1 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_1 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_1 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_1 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_1 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_1 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_1 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_1 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_1 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_1 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_1 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_1 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_1 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_1 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_1 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_1 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_1 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_1 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_1 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_1 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_1 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_1 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_1 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_1 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_1 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_1 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_1 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_1 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_1 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_1 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_1 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_1 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_1 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_1 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_1 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_1 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_1 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_1 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_1 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_1 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_1 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_1 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_1 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_1 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_1 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_1 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_1 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_1 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_1 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_1 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_1 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_1 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_1 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_1 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_1 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_1 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_1 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_1 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_1 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_1 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_1 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_1 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_1_3)
      8'b00000000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_1_2 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_1_2 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_1_5)
      8'b00000000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_1_4 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_1_4 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(_zz__zz_roundKeyReg_0_1_7)
      8'b00000000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_0;
      8'b00000001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_1;
      8'b00000010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_2;
      8'b00000011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_3;
      8'b00000100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_4;
      8'b00000101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_5;
      8'b00000110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_6;
      8'b00000111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_7;
      8'b00001000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_8;
      8'b00001001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_9;
      8'b00001010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_10;
      8'b00001011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_11;
      8'b00001100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_12;
      8'b00001101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_13;
      8'b00001110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_14;
      8'b00001111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_15;
      8'b00010000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_16;
      8'b00010001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_17;
      8'b00010010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_18;
      8'b00010011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_19;
      8'b00010100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_20;
      8'b00010101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_21;
      8'b00010110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_22;
      8'b00010111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_23;
      8'b00011000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_24;
      8'b00011001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_25;
      8'b00011010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_26;
      8'b00011011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_27;
      8'b00011100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_28;
      8'b00011101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_29;
      8'b00011110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_30;
      8'b00011111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_31;
      8'b00100000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_32;
      8'b00100001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_33;
      8'b00100010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_34;
      8'b00100011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_35;
      8'b00100100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_36;
      8'b00100101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_37;
      8'b00100110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_38;
      8'b00100111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_39;
      8'b00101000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_40;
      8'b00101001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_41;
      8'b00101010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_42;
      8'b00101011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_43;
      8'b00101100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_44;
      8'b00101101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_45;
      8'b00101110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_46;
      8'b00101111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_47;
      8'b00110000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_48;
      8'b00110001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_49;
      8'b00110010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_50;
      8'b00110011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_51;
      8'b00110100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_52;
      8'b00110101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_53;
      8'b00110110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_54;
      8'b00110111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_55;
      8'b00111000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_56;
      8'b00111001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_57;
      8'b00111010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_58;
      8'b00111011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_59;
      8'b00111100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_60;
      8'b00111101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_61;
      8'b00111110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_62;
      8'b00111111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_63;
      8'b01000000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_64;
      8'b01000001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_65;
      8'b01000010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_66;
      8'b01000011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_67;
      8'b01000100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_68;
      8'b01000101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_69;
      8'b01000110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_70;
      8'b01000111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_71;
      8'b01001000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_72;
      8'b01001001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_73;
      8'b01001010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_74;
      8'b01001011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_75;
      8'b01001100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_76;
      8'b01001101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_77;
      8'b01001110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_78;
      8'b01001111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_79;
      8'b01010000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_80;
      8'b01010001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_81;
      8'b01010010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_82;
      8'b01010011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_83;
      8'b01010100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_84;
      8'b01010101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_85;
      8'b01010110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_86;
      8'b01010111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_87;
      8'b01011000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_88;
      8'b01011001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_89;
      8'b01011010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_90;
      8'b01011011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_91;
      8'b01011100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_92;
      8'b01011101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_93;
      8'b01011110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_94;
      8'b01011111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_95;
      8'b01100000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_96;
      8'b01100001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_97;
      8'b01100010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_98;
      8'b01100011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_99;
      8'b01100100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_100;
      8'b01100101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_101;
      8'b01100110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_102;
      8'b01100111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_103;
      8'b01101000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_104;
      8'b01101001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_105;
      8'b01101010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_106;
      8'b01101011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_107;
      8'b01101100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_108;
      8'b01101101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_109;
      8'b01101110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_110;
      8'b01101111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_111;
      8'b01110000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_112;
      8'b01110001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_113;
      8'b01110010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_114;
      8'b01110011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_115;
      8'b01110100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_116;
      8'b01110101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_117;
      8'b01110110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_118;
      8'b01110111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_119;
      8'b01111000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_120;
      8'b01111001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_121;
      8'b01111010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_122;
      8'b01111011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_123;
      8'b01111100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_124;
      8'b01111101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_125;
      8'b01111110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_126;
      8'b01111111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_127;
      8'b10000000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_128;
      8'b10000001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_129;
      8'b10000010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_130;
      8'b10000011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_131;
      8'b10000100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_132;
      8'b10000101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_133;
      8'b10000110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_134;
      8'b10000111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_135;
      8'b10001000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_136;
      8'b10001001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_137;
      8'b10001010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_138;
      8'b10001011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_139;
      8'b10001100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_140;
      8'b10001101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_141;
      8'b10001110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_142;
      8'b10001111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_143;
      8'b10010000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_144;
      8'b10010001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_145;
      8'b10010010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_146;
      8'b10010011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_147;
      8'b10010100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_148;
      8'b10010101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_149;
      8'b10010110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_150;
      8'b10010111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_151;
      8'b10011000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_152;
      8'b10011001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_153;
      8'b10011010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_154;
      8'b10011011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_155;
      8'b10011100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_156;
      8'b10011101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_157;
      8'b10011110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_158;
      8'b10011111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_159;
      8'b10100000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_160;
      8'b10100001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_161;
      8'b10100010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_162;
      8'b10100011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_163;
      8'b10100100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_164;
      8'b10100101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_165;
      8'b10100110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_166;
      8'b10100111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_167;
      8'b10101000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_168;
      8'b10101001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_169;
      8'b10101010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_170;
      8'b10101011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_171;
      8'b10101100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_172;
      8'b10101101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_173;
      8'b10101110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_174;
      8'b10101111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_175;
      8'b10110000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_176;
      8'b10110001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_177;
      8'b10110010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_178;
      8'b10110011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_179;
      8'b10110100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_180;
      8'b10110101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_181;
      8'b10110110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_182;
      8'b10110111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_183;
      8'b10111000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_184;
      8'b10111001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_185;
      8'b10111010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_186;
      8'b10111011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_187;
      8'b10111100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_188;
      8'b10111101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_189;
      8'b10111110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_190;
      8'b10111111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_191;
      8'b11000000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_192;
      8'b11000001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_193;
      8'b11000010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_194;
      8'b11000011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_195;
      8'b11000100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_196;
      8'b11000101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_197;
      8'b11000110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_198;
      8'b11000111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_199;
      8'b11001000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_200;
      8'b11001001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_201;
      8'b11001010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_202;
      8'b11001011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_203;
      8'b11001100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_204;
      8'b11001101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_205;
      8'b11001110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_206;
      8'b11001111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_207;
      8'b11010000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_208;
      8'b11010001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_209;
      8'b11010010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_210;
      8'b11010011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_211;
      8'b11010100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_212;
      8'b11010101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_213;
      8'b11010110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_214;
      8'b11010111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_215;
      8'b11011000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_216;
      8'b11011001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_217;
      8'b11011010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_218;
      8'b11011011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_219;
      8'b11011100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_220;
      8'b11011101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_221;
      8'b11011110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_222;
      8'b11011111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_223;
      8'b11100000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_224;
      8'b11100001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_225;
      8'b11100010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_226;
      8'b11100011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_227;
      8'b11100100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_228;
      8'b11100101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_229;
      8'b11100110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_230;
      8'b11100111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_231;
      8'b11101000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_232;
      8'b11101001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_233;
      8'b11101010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_234;
      8'b11101011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_235;
      8'b11101100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_236;
      8'b11101101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_237;
      8'b11101110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_238;
      8'b11101111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_239;
      8'b11110000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_240;
      8'b11110001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_241;
      8'b11110010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_242;
      8'b11110011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_243;
      8'b11110100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_244;
      8'b11110101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_245;
      8'b11110110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_246;
      8'b11110111 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_247;
      8'b11111000 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_248;
      8'b11111001 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_249;
      8'b11111010 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_250;
      8'b11111011 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_251;
      8'b11111100 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_252;
      8'b11111101 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_253;
      8'b11111110 : _zz__zz_roundKeyReg_0_1_6 = sboxRom_254;
      default : _zz__zz_roundKeyReg_0_1_6 = sboxRom_255;
    endcase
  end

  always @(*) begin
    case(rconCounter)
      4'b0000 : _zz__zz_roundKeyReg_0_1_8 = rcon_0;
      4'b0001 : _zz__zz_roundKeyReg_0_1_8 = rcon_1;
      4'b0010 : _zz__zz_roundKeyReg_0_1_8 = rcon_2;
      4'b0011 : _zz__zz_roundKeyReg_0_1_8 = rcon_3;
      4'b0100 : _zz__zz_roundKeyReg_0_1_8 = rcon_4;
      4'b0101 : _zz__zz_roundKeyReg_0_1_8 = rcon_5;
      4'b0110 : _zz__zz_roundKeyReg_0_1_8 = rcon_6;
      4'b0111 : _zz__zz_roundKeyReg_0_1_8 = rcon_7;
      4'b1000 : _zz__zz_roundKeyReg_0_1_8 = rcon_8;
      default : _zz__zz_roundKeyReg_0_1_8 = rcon_9;
    endcase
  end

  assign sboxRom_0 = 8'h63;
  assign sboxRom_1 = 8'h7c;
  assign sboxRom_2 = 8'h77;
  assign sboxRom_3 = 8'h7b;
  assign sboxRom_4 = 8'hf2;
  assign sboxRom_5 = 8'h6b;
  assign sboxRom_6 = 8'h6f;
  assign sboxRom_7 = 8'hc5;
  assign sboxRom_8 = 8'h30;
  assign sboxRom_9 = 8'h01;
  assign sboxRom_10 = 8'h67;
  assign sboxRom_11 = 8'h2b;
  assign sboxRom_12 = 8'hfe;
  assign sboxRom_13 = 8'hd7;
  assign sboxRom_14 = 8'hab;
  assign sboxRom_15 = 8'h76;
  assign sboxRom_16 = 8'hca;
  assign sboxRom_17 = 8'h82;
  assign sboxRom_18 = 8'hc9;
  assign sboxRom_19 = 8'h7d;
  assign sboxRom_20 = 8'hfa;
  assign sboxRom_21 = 8'h59;
  assign sboxRom_22 = 8'h47;
  assign sboxRom_23 = 8'hf0;
  assign sboxRom_24 = 8'had;
  assign sboxRom_25 = 8'hd4;
  assign sboxRom_26 = 8'ha2;
  assign sboxRom_27 = 8'haf;
  assign sboxRom_28 = 8'h9c;
  assign sboxRom_29 = 8'ha4;
  assign sboxRom_30 = 8'h72;
  assign sboxRom_31 = 8'hc0;
  assign sboxRom_32 = 8'hb7;
  assign sboxRom_33 = 8'hfd;
  assign sboxRom_34 = 8'h93;
  assign sboxRom_35 = 8'h26;
  assign sboxRom_36 = 8'h36;
  assign sboxRom_37 = 8'h3f;
  assign sboxRom_38 = 8'hf7;
  assign sboxRom_39 = 8'hcc;
  assign sboxRom_40 = 8'h34;
  assign sboxRom_41 = 8'ha5;
  assign sboxRom_42 = 8'he5;
  assign sboxRom_43 = 8'hf1;
  assign sboxRom_44 = 8'h71;
  assign sboxRom_45 = 8'hd8;
  assign sboxRom_46 = 8'h31;
  assign sboxRom_47 = 8'h15;
  assign sboxRom_48 = 8'h04;
  assign sboxRom_49 = 8'hc7;
  assign sboxRom_50 = 8'h23;
  assign sboxRom_51 = 8'hc3;
  assign sboxRom_52 = 8'h18;
  assign sboxRom_53 = 8'h96;
  assign sboxRom_54 = 8'h05;
  assign sboxRom_55 = 8'h9a;
  assign sboxRom_56 = 8'h07;
  assign sboxRom_57 = 8'h12;
  assign sboxRom_58 = 8'h80;
  assign sboxRom_59 = 8'he2;
  assign sboxRom_60 = 8'heb;
  assign sboxRom_61 = 8'h27;
  assign sboxRom_62 = 8'hb2;
  assign sboxRom_63 = 8'h75;
  assign sboxRom_64 = 8'h09;
  assign sboxRom_65 = 8'h83;
  assign sboxRom_66 = 8'h2c;
  assign sboxRom_67 = 8'h1a;
  assign sboxRom_68 = 8'h1b;
  assign sboxRom_69 = 8'h6e;
  assign sboxRom_70 = 8'h5a;
  assign sboxRom_71 = 8'ha0;
  assign sboxRom_72 = 8'h52;
  assign sboxRom_73 = 8'h3b;
  assign sboxRom_74 = 8'hd6;
  assign sboxRom_75 = 8'hb3;
  assign sboxRom_76 = 8'h29;
  assign sboxRom_77 = 8'he3;
  assign sboxRom_78 = 8'h2f;
  assign sboxRom_79 = 8'h84;
  assign sboxRom_80 = 8'h53;
  assign sboxRom_81 = 8'hd1;
  assign sboxRom_82 = 8'h0;
  assign sboxRom_83 = 8'hed;
  assign sboxRom_84 = 8'h20;
  assign sboxRom_85 = 8'hfc;
  assign sboxRom_86 = 8'hb1;
  assign sboxRom_87 = 8'h5b;
  assign sboxRom_88 = 8'h6a;
  assign sboxRom_89 = 8'hcb;
  assign sboxRom_90 = 8'hbe;
  assign sboxRom_91 = 8'h39;
  assign sboxRom_92 = 8'h4a;
  assign sboxRom_93 = 8'h4c;
  assign sboxRom_94 = 8'h58;
  assign sboxRom_95 = 8'hcf;
  assign sboxRom_96 = 8'hd0;
  assign sboxRom_97 = 8'hef;
  assign sboxRom_98 = 8'haa;
  assign sboxRom_99 = 8'hfb;
  assign sboxRom_100 = 8'h43;
  assign sboxRom_101 = 8'h4d;
  assign sboxRom_102 = 8'h33;
  assign sboxRom_103 = 8'h85;
  assign sboxRom_104 = 8'h45;
  assign sboxRom_105 = 8'hf9;
  assign sboxRom_106 = 8'h02;
  assign sboxRom_107 = 8'h7f;
  assign sboxRom_108 = 8'h50;
  assign sboxRom_109 = 8'h3c;
  assign sboxRom_110 = 8'h9f;
  assign sboxRom_111 = 8'ha8;
  assign sboxRom_112 = 8'h51;
  assign sboxRom_113 = 8'ha3;
  assign sboxRom_114 = 8'h40;
  assign sboxRom_115 = 8'h8f;
  assign sboxRom_116 = 8'h92;
  assign sboxRom_117 = 8'h9d;
  assign sboxRom_118 = 8'h38;
  assign sboxRom_119 = 8'hf5;
  assign sboxRom_120 = 8'hbc;
  assign sboxRom_121 = 8'hb6;
  assign sboxRom_122 = 8'hda;
  assign sboxRom_123 = 8'h21;
  assign sboxRom_124 = 8'h10;
  assign sboxRom_125 = 8'hff;
  assign sboxRom_126 = 8'hf3;
  assign sboxRom_127 = 8'hd2;
  assign sboxRom_128 = 8'hcd;
  assign sboxRom_129 = 8'h0c;
  assign sboxRom_130 = 8'h13;
  assign sboxRom_131 = 8'hec;
  assign sboxRom_132 = 8'h5f;
  assign sboxRom_133 = 8'h97;
  assign sboxRom_134 = 8'h44;
  assign sboxRom_135 = 8'h17;
  assign sboxRom_136 = 8'hc4;
  assign sboxRom_137 = 8'ha7;
  assign sboxRom_138 = 8'h7e;
  assign sboxRom_139 = 8'h3d;
  assign sboxRom_140 = 8'h64;
  assign sboxRom_141 = 8'h5d;
  assign sboxRom_142 = 8'h19;
  assign sboxRom_143 = 8'h73;
  assign sboxRom_144 = 8'h60;
  assign sboxRom_145 = 8'h81;
  assign sboxRom_146 = 8'h4f;
  assign sboxRom_147 = 8'hdc;
  assign sboxRom_148 = 8'h22;
  assign sboxRom_149 = 8'h2a;
  assign sboxRom_150 = 8'h90;
  assign sboxRom_151 = 8'h88;
  assign sboxRom_152 = 8'h46;
  assign sboxRom_153 = 8'hee;
  assign sboxRom_154 = 8'hb8;
  assign sboxRom_155 = 8'h14;
  assign sboxRom_156 = 8'hde;
  assign sboxRom_157 = 8'h5e;
  assign sboxRom_158 = 8'h0b;
  assign sboxRom_159 = 8'hdb;
  assign sboxRom_160 = 8'he0;
  assign sboxRom_161 = 8'h32;
  assign sboxRom_162 = 8'h3a;
  assign sboxRom_163 = 8'h0a;
  assign sboxRom_164 = 8'h49;
  assign sboxRom_165 = 8'h06;
  assign sboxRom_166 = 8'h24;
  assign sboxRom_167 = 8'h5c;
  assign sboxRom_168 = 8'hc2;
  assign sboxRom_169 = 8'hd3;
  assign sboxRom_170 = 8'hac;
  assign sboxRom_171 = 8'h62;
  assign sboxRom_172 = 8'h91;
  assign sboxRom_173 = 8'h95;
  assign sboxRom_174 = 8'he4;
  assign sboxRom_175 = 8'h79;
  assign sboxRom_176 = 8'he7;
  assign sboxRom_177 = 8'hc8;
  assign sboxRom_178 = 8'h37;
  assign sboxRom_179 = 8'h6d;
  assign sboxRom_180 = 8'h8d;
  assign sboxRom_181 = 8'hd5;
  assign sboxRom_182 = 8'h4e;
  assign sboxRom_183 = 8'ha9;
  assign sboxRom_184 = 8'h6c;
  assign sboxRom_185 = 8'h56;
  assign sboxRom_186 = 8'hf4;
  assign sboxRom_187 = 8'hea;
  assign sboxRom_188 = 8'h65;
  assign sboxRom_189 = 8'h7a;
  assign sboxRom_190 = 8'hae;
  assign sboxRom_191 = 8'h08;
  assign sboxRom_192 = 8'hba;
  assign sboxRom_193 = 8'h78;
  assign sboxRom_194 = 8'h25;
  assign sboxRom_195 = 8'h2e;
  assign sboxRom_196 = 8'h1c;
  assign sboxRom_197 = 8'ha6;
  assign sboxRom_198 = 8'hb4;
  assign sboxRom_199 = 8'hc6;
  assign sboxRom_200 = 8'he8;
  assign sboxRom_201 = 8'hdd;
  assign sboxRom_202 = 8'h74;
  assign sboxRom_203 = 8'h1f;
  assign sboxRom_204 = 8'h4b;
  assign sboxRom_205 = 8'hbd;
  assign sboxRom_206 = 8'h8b;
  assign sboxRom_207 = 8'h8a;
  assign sboxRom_208 = 8'h70;
  assign sboxRom_209 = 8'h3e;
  assign sboxRom_210 = 8'hb5;
  assign sboxRom_211 = 8'h66;
  assign sboxRom_212 = 8'h48;
  assign sboxRom_213 = 8'h03;
  assign sboxRom_214 = 8'hf6;
  assign sboxRom_215 = 8'h0e;
  assign sboxRom_216 = 8'h61;
  assign sboxRom_217 = 8'h35;
  assign sboxRom_218 = 8'h57;
  assign sboxRom_219 = 8'hb9;
  assign sboxRom_220 = 8'h86;
  assign sboxRom_221 = 8'hc1;
  assign sboxRom_222 = 8'h1d;
  assign sboxRom_223 = 8'h9e;
  assign sboxRom_224 = 8'he1;
  assign sboxRom_225 = 8'hf8;
  assign sboxRom_226 = 8'h98;
  assign sboxRom_227 = 8'h11;
  assign sboxRom_228 = 8'h69;
  assign sboxRom_229 = 8'hd9;
  assign sboxRom_230 = 8'h8e;
  assign sboxRom_231 = 8'h94;
  assign sboxRom_232 = 8'h9b;
  assign sboxRom_233 = 8'h1e;
  assign sboxRom_234 = 8'h87;
  assign sboxRom_235 = 8'he9;
  assign sboxRom_236 = 8'hce;
  assign sboxRom_237 = 8'h55;
  assign sboxRom_238 = 8'h28;
  assign sboxRom_239 = 8'hdf;
  assign sboxRom_240 = 8'h8c;
  assign sboxRom_241 = 8'ha1;
  assign sboxRom_242 = 8'h89;
  assign sboxRom_243 = 8'h0d;
  assign sboxRom_244 = 8'hbf;
  assign sboxRom_245 = 8'he6;
  assign sboxRom_246 = 8'h42;
  assign sboxRom_247 = 8'h68;
  assign sboxRom_248 = 8'h41;
  assign sboxRom_249 = 8'h99;
  assign sboxRom_250 = 8'h2d;
  assign sboxRom_251 = 8'h0f;
  assign sboxRom_252 = 8'hb0;
  assign sboxRom_253 = 8'h54;
  assign sboxRom_254 = 8'hbb;
  assign sboxRom_255 = 8'h16;
  assign rcon_0 = 8'h01;
  assign rcon_1 = 8'h02;
  assign rcon_2 = 8'h04;
  assign rcon_3 = 8'h08;
  assign rcon_4 = 8'h10;
  assign rcon_5 = 8'h20;
  assign rcon_6 = 8'h40;
  assign rcon_7 = 8'h80;
  assign rcon_8 = 8'h1b;
  assign rcon_9 = 8'h36;
  assign io_busy = running;
  always @(*) begin
    io_done = 1'b0;
    if(!when_AES128_l150) begin
      if(running) begin
        if(when_AES128_l227) begin
          io_done = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_dataOut = stateReg;
    if(!when_AES128_l150) begin
      if(running) begin
        if(when_AES128_l227) begin
          io_dataOut = stateReg;
        end
      end
    end
  end

  always @(*) begin
    newStateComb = 128'h0;
    if(!when_AES128_l150) begin
      if(running) begin
        newStateComb = _zz_stateReg_68;
      end
    end
  end

  always @(*) begin
    rkBitsUsedComb = 128'h0;
    if(!when_AES128_l150) begin
      if(running) begin
        rkBitsUsedComb = _zz_stateReg_69;
      end
    end
  end

  assign when_AES128_l150 = (io_start && (! running));
  assign _zz_stateReg = io_key[127 : 96];
  assign _zz_stateReg_1 = io_key[95 : 64];
  assign _zz_stateReg_2 = io_key[63 : 32];
  assign _zz_stateReg_3 = io_key[31 : 0];
  assign _zz_stateReg_4 = _zz__zz_stateReg_4;
  assign _zz_stateReg_8 = _zz__zz_stateReg_8;
  assign _zz_stateReg_12 = _zz__zz_stateReg_12;
  assign _zz_stateReg_16 = _zz__zz_stateReg_16;
  assign _zz_stateReg_5 = _zz__zz_stateReg_5;
  assign _zz_stateReg_9 = _zz__zz_stateReg_9;
  assign _zz_stateReg_13 = _zz__zz_stateReg_13;
  assign _zz_stateReg_17 = _zz__zz_stateReg_17;
  assign _zz_stateReg_6 = _zz__zz_stateReg_6;
  assign _zz_stateReg_10 = _zz__zz_stateReg_10;
  assign _zz_stateReg_14 = _zz__zz_stateReg_14;
  assign _zz_stateReg_18 = _zz__zz_stateReg_18;
  assign _zz_stateReg_7 = _zz__zz_stateReg_7;
  assign _zz_stateReg_11 = _zz__zz_stateReg_11;
  assign _zz_stateReg_15 = _zz__zz_stateReg_15;
  assign _zz_stateReg_19 = _zz__zz_stateReg_19;
  assign when_AES128_l192 = (roundCount == 4'b1001);
  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_20 = _zz_stateReg_4;
    end else begin
      _zz_stateReg_20 = ((((_zz_stateReg_4[7] ? (_zz_stateReg_36 ^ 8'h1b) : _zz_stateReg_36) ^ ((_zz_stateReg_5[7] ? (_zz_stateReg_37 ^ 8'h1b) : _zz_stateReg_37) ^ _zz_stateReg_5)) ^ _zz_stateReg_6) ^ _zz_stateReg_7);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_21 = _zz_stateReg_5;
    end else begin
      _zz_stateReg_21 = (((_zz_stateReg_4 ^ (_zz_stateReg_5[7] ? (_zz_stateReg_38 ^ 8'h1b) : _zz_stateReg_38)) ^ ((_zz_stateReg_6[7] ? (_zz_stateReg_39 ^ 8'h1b) : _zz_stateReg_39) ^ _zz_stateReg_6)) ^ _zz_stateReg_7);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_22 = _zz_stateReg_6;
    end else begin
      _zz_stateReg_22 = (((_zz_stateReg_4 ^ _zz_stateReg_5) ^ (_zz_stateReg_6[7] ? (_zz_stateReg_40 ^ 8'h1b) : _zz_stateReg_40)) ^ ((_zz_stateReg_7[7] ? (_zz_stateReg_41 ^ 8'h1b) : _zz_stateReg_41) ^ _zz_stateReg_7));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_23 = _zz_stateReg_7;
    end else begin
      _zz_stateReg_23 = (((((_zz_stateReg_4[7] ? (_zz_stateReg_42 ^ 8'h1b) : _zz_stateReg_42) ^ _zz_stateReg_4) ^ _zz_stateReg_5) ^ _zz_stateReg_6) ^ (_zz_stateReg_7[7] ? (_zz_stateReg_43 ^ 8'h1b) : _zz_stateReg_43));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_24 = _zz_stateReg_8;
    end else begin
      _zz_stateReg_24 = ((((_zz_stateReg_8[7] ? (_zz_stateReg_44 ^ 8'h1b) : _zz_stateReg_44) ^ ((_zz_stateReg_9[7] ? (_zz_stateReg_45 ^ 8'h1b) : _zz_stateReg_45) ^ _zz_stateReg_9)) ^ _zz_stateReg_10) ^ _zz_stateReg_11);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_25 = _zz_stateReg_9;
    end else begin
      _zz_stateReg_25 = (((_zz_stateReg_8 ^ (_zz_stateReg_9[7] ? (_zz_stateReg_46 ^ 8'h1b) : _zz_stateReg_46)) ^ ((_zz_stateReg_10[7] ? (_zz_stateReg_47 ^ 8'h1b) : _zz_stateReg_47) ^ _zz_stateReg_10)) ^ _zz_stateReg_11);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_26 = _zz_stateReg_10;
    end else begin
      _zz_stateReg_26 = (((_zz_stateReg_8 ^ _zz_stateReg_9) ^ (_zz_stateReg_10[7] ? (_zz_stateReg_48 ^ 8'h1b) : _zz_stateReg_48)) ^ ((_zz_stateReg_11[7] ? (_zz_stateReg_49 ^ 8'h1b) : _zz_stateReg_49) ^ _zz_stateReg_11));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_27 = _zz_stateReg_11;
    end else begin
      _zz_stateReg_27 = (((((_zz_stateReg_8[7] ? (_zz_stateReg_50 ^ 8'h1b) : _zz_stateReg_50) ^ _zz_stateReg_8) ^ _zz_stateReg_9) ^ _zz_stateReg_10) ^ (_zz_stateReg_11[7] ? (_zz_stateReg_51 ^ 8'h1b) : _zz_stateReg_51));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_28 = _zz_stateReg_12;
    end else begin
      _zz_stateReg_28 = ((((_zz_stateReg_12[7] ? (_zz_stateReg_52 ^ 8'h1b) : _zz_stateReg_52) ^ ((_zz_stateReg_13[7] ? (_zz_stateReg_53 ^ 8'h1b) : _zz_stateReg_53) ^ _zz_stateReg_13)) ^ _zz_stateReg_14) ^ _zz_stateReg_15);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_29 = _zz_stateReg_13;
    end else begin
      _zz_stateReg_29 = (((_zz_stateReg_12 ^ (_zz_stateReg_13[7] ? (_zz_stateReg_54 ^ 8'h1b) : _zz_stateReg_54)) ^ ((_zz_stateReg_14[7] ? (_zz_stateReg_55 ^ 8'h1b) : _zz_stateReg_55) ^ _zz_stateReg_14)) ^ _zz_stateReg_15);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_30 = _zz_stateReg_14;
    end else begin
      _zz_stateReg_30 = (((_zz_stateReg_12 ^ _zz_stateReg_13) ^ (_zz_stateReg_14[7] ? (_zz_stateReg_56 ^ 8'h1b) : _zz_stateReg_56)) ^ ((_zz_stateReg_15[7] ? (_zz_stateReg_57 ^ 8'h1b) : _zz_stateReg_57) ^ _zz_stateReg_15));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_31 = _zz_stateReg_15;
    end else begin
      _zz_stateReg_31 = (((((_zz_stateReg_12[7] ? (_zz_stateReg_58 ^ 8'h1b) : _zz_stateReg_58) ^ _zz_stateReg_12) ^ _zz_stateReg_13) ^ _zz_stateReg_14) ^ (_zz_stateReg_15[7] ? (_zz_stateReg_59 ^ 8'h1b) : _zz_stateReg_59));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_32 = _zz_stateReg_16;
    end else begin
      _zz_stateReg_32 = ((((_zz_stateReg_16[7] ? (_zz_stateReg_60 ^ 8'h1b) : _zz_stateReg_60) ^ ((_zz_stateReg_17[7] ? (_zz_stateReg_61 ^ 8'h1b) : _zz_stateReg_61) ^ _zz_stateReg_17)) ^ _zz_stateReg_18) ^ _zz_stateReg_19);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_33 = _zz_stateReg_17;
    end else begin
      _zz_stateReg_33 = (((_zz_stateReg_16 ^ (_zz_stateReg_17[7] ? (_zz_stateReg_62 ^ 8'h1b) : _zz_stateReg_62)) ^ ((_zz_stateReg_18[7] ? (_zz_stateReg_63 ^ 8'h1b) : _zz_stateReg_63) ^ _zz_stateReg_18)) ^ _zz_stateReg_19);
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_34 = _zz_stateReg_18;
    end else begin
      _zz_stateReg_34 = (((_zz_stateReg_16 ^ _zz_stateReg_17) ^ (_zz_stateReg_18[7] ? (_zz_stateReg_64 ^ 8'h1b) : _zz_stateReg_64)) ^ ((_zz_stateReg_19[7] ? (_zz_stateReg_65 ^ 8'h1b) : _zz_stateReg_65) ^ _zz_stateReg_19));
    end
  end

  always @(*) begin
    if(when_AES128_l192) begin
      _zz_stateReg_35 = _zz_stateReg_19;
    end else begin
      _zz_stateReg_35 = (((((_zz_stateReg_16[7] ? (_zz_stateReg_66 ^ 8'h1b) : _zz_stateReg_66) ^ _zz_stateReg_16) ^ _zz_stateReg_17) ^ _zz_stateReg_18) ^ (_zz_stateReg_19[7] ? (_zz_stateReg_67 ^ 8'h1b) : _zz_stateReg_67));
    end
  end

  assign _zz_stateReg_36 = _zz__zz_stateReg_36[7 : 0];
  assign _zz_stateReg_37 = _zz__zz_stateReg_37[7 : 0];
  assign _zz_stateReg_38 = _zz__zz_stateReg_38[7 : 0];
  assign _zz_stateReg_39 = _zz__zz_stateReg_39[7 : 0];
  assign _zz_stateReg_40 = _zz__zz_stateReg_40[7 : 0];
  assign _zz_stateReg_41 = _zz__zz_stateReg_41[7 : 0];
  assign _zz_stateReg_42 = _zz__zz_stateReg_42[7 : 0];
  assign _zz_stateReg_43 = _zz__zz_stateReg_43[7 : 0];
  assign _zz_stateReg_44 = _zz__zz_stateReg_44[7 : 0];
  assign _zz_stateReg_45 = _zz__zz_stateReg_45[7 : 0];
  assign _zz_stateReg_46 = _zz__zz_stateReg_46[7 : 0];
  assign _zz_stateReg_47 = _zz__zz_stateReg_47[7 : 0];
  assign _zz_stateReg_48 = _zz__zz_stateReg_48[7 : 0];
  assign _zz_stateReg_49 = _zz__zz_stateReg_49[7 : 0];
  assign _zz_stateReg_50 = _zz__zz_stateReg_50[7 : 0];
  assign _zz_stateReg_51 = _zz__zz_stateReg_51[7 : 0];
  assign _zz_stateReg_52 = _zz__zz_stateReg_52[7 : 0];
  assign _zz_stateReg_53 = _zz__zz_stateReg_53[7 : 0];
  assign _zz_stateReg_54 = _zz__zz_stateReg_54[7 : 0];
  assign _zz_stateReg_55 = _zz__zz_stateReg_55[7 : 0];
  assign _zz_stateReg_56 = _zz__zz_stateReg_56[7 : 0];
  assign _zz_stateReg_57 = _zz__zz_stateReg_57[7 : 0];
  assign _zz_stateReg_58 = _zz__zz_stateReg_58[7 : 0];
  assign _zz_stateReg_59 = _zz__zz_stateReg_59[7 : 0];
  assign _zz_stateReg_60 = _zz__zz_stateReg_60[7 : 0];
  assign _zz_stateReg_61 = _zz__zz_stateReg_61[7 : 0];
  assign _zz_stateReg_62 = _zz__zz_stateReg_62[7 : 0];
  assign _zz_stateReg_63 = _zz__zz_stateReg_63[7 : 0];
  assign _zz_stateReg_64 = _zz__zz_stateReg_64[7 : 0];
  assign _zz_stateReg_65 = _zz__zz_stateReg_65[7 : 0];
  assign _zz_stateReg_66 = _zz__zz_stateReg_66[7 : 0];
  assign _zz_stateReg_67 = _zz__zz_stateReg_67[7 : 0];
  assign _zz_stateReg_68 = {{{{{{{{{{{_zz__zz_stateReg_68,_zz__zz_stateReg_68_1},_zz_stateReg_26},_zz_stateReg_27},_zz_stateReg_28},_zz_stateReg_29},_zz_stateReg_30},_zz_stateReg_31},_zz_stateReg_32},_zz_stateReg_33},_zz_stateReg_34},_zz_stateReg_35};
  assign _zz_roundKeyReg_0 = {roundKeyReg_3[23 : 0],roundKeyReg_3[31 : 24]};
  assign _zz_roundKeyReg_0_1 = (roundKeyReg_0 ^ ({{{_zz__zz_roundKeyReg_0_1,_zz__zz_roundKeyReg_0_1_2},_zz__zz_roundKeyReg_0_1_4},_zz__zz_roundKeyReg_0_1_6} ^ {_zz__zz_roundKeyReg_0_1_8,24'h0}));
  assign _zz_roundKeyReg_1 = (roundKeyReg_1 ^ _zz_roundKeyReg_0_1);
  assign _zz_roundKeyReg_2 = (roundKeyReg_2 ^ _zz_roundKeyReg_1);
  assign _zz_roundKeyReg_3 = (roundKeyReg_3 ^ _zz_roundKeyReg_2);
  assign _zz_stateReg_69 = {{{{{{{{{_zz__zz_stateReg_69,_zz__zz_stateReg_69_1},_zz__zz_stateReg_69_2},_zz_roundKeyReg_2[23 : 16]},_zz_roundKeyReg_2[15 : 8]},_zz_roundKeyReg_2[7 : 0]},_zz_roundKeyReg_3[31 : 24]},_zz_roundKeyReg_3[23 : 16]},_zz_roundKeyReg_3[15 : 8]},_zz_roundKeyReg_3[7 : 0]};
  assign when_AES128_l227 = (roundCount == 4'b1010);
  assign when_AES128_l233 = (rconCounter < 4'b1001);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      stateReg <= 128'h0;
      roundKeyReg_0 <= 32'h0;
      roundKeyReg_1 <= 32'h0;
      roundKeyReg_2 <= 32'h0;
      roundKeyReg_3 <= 32'h0;
      roundCount <= 4'b0000;
      running <= 1'b0;
      rconCounter <= 4'b0000;
    end else begin
      if(when_AES128_l150) begin
        running <= 1'b1;
        stateReg <= {{{{{{_zz_stateReg_70,_zz_stateReg_82},_zz_stateReg_83},(_zz_stateReg_84 ^ _zz_stateReg_85)},(_zz_stateReg_86 ^ _zz_stateReg_3[23 : 16])},(io_dataIn[15 : 8] ^ _zz_stateReg_3[15 : 8])},(io_dataIn[7 : 0] ^ _zz_stateReg_3[7 : 0])};
        roundKeyReg_0 <= _zz_stateReg;
        roundKeyReg_1 <= _zz_stateReg_1;
        roundKeyReg_2 <= _zz_stateReg_2;
        roundKeyReg_3 <= _zz_stateReg_3;
        roundCount <= 4'b0000;
        rconCounter <= 4'b0000;
      end else begin
        if(running) begin
          stateReg <= (_zz_stateReg_68 ^ _zz_stateReg_69);
          roundKeyReg_0 <= _zz_roundKeyReg_0_1;
          roundKeyReg_1 <= _zz_roundKeyReg_1;
          roundKeyReg_2 <= _zz_roundKeyReg_2;
          roundKeyReg_3 <= _zz_roundKeyReg_3;
          if(when_AES128_l227) begin
            running <= 1'b0;
          end else begin
            roundCount <= (roundCount + 4'b0001);
            if(when_AES128_l233) begin
              rconCounter <= (rconCounter + 4'b0001);
            end
          end
        end
      end
    end
  end


endmodule
